module IFU(
  input          clock,
  input          reset,
  output         io_imem_valid,
  output [31:0]  io_imem_addr,
  output         io_imem_fence,
  input          io_imem_fence_finish,
  input          io_imem_data_ok,
  input  [127:0] io_imem_inst,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_pc,
  output [127:0] io_out_bits_inst,
  output         io_out_bits_uncache,
  output [1:0]   io_out_bits_offset,
  output [1:0]   io_out_bits_bp_br_offset,
  output         io_out_bits_bp_br_taken,
  output [31:0]  io_out_bits_bp_br_target,
  output [1:0]   io_out_bits_bp_br_type,
  input          io_reflush_bus_is_reflush,
  input  [31:0]  io_reflush_bus_br_target,
  output         io_bpu_valid,
  output [31:0]  io_bpu_pc,
  input          io_bpu_bp_ok,
  input          io_bpu_bp_taken,
  input  [31:0]  io_bpu_bp_target,
  input  [1:0]   io_bpu_bp_offset,
  output         io_bpu_is_reflush,
  input  [1:0]   io_bpu_bp_type,
  output [2:0]   io_bpu_call_count,
  output [2:0]   io_bpu_ret_count,
  input          dcache_fence_finish_0,
  input          fence_i,
  output         icache_fence_finish_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] pc; // @[IFU.scala 14:19]
  reg [31:0] bp_pc_reg; // @[IFU.scala 16:26]
  reg  bp_taken_reg; // @[IFU.scala 18:29]
  reg [1:0] bp_type_reg; // @[IFU.scala 20:28]
  reg [1:0] bp_offset_reg; // @[IFU.scala 22:30]
  reg [31:0] bpu_reg_pc; // @[IFU.scala 24:27]
  reg  imem_reg_valid; // @[IFU.scala 25:31]
  wire  bp_taken = io_bpu_bp_ok ? io_bpu_bp_taken : bp_taken_reg; // @[IFU.scala 40:18]
  wire [31:0] bp_pc = io_bpu_bp_ok ? io_bpu_bp_target : bp_pc_reg; // @[IFU.scala 41:15]
  wire [1:0] bp_type = io_bpu_bp_ok ? io_bpu_bp_type : bp_type_reg; // @[IFU.scala 42:17]
  reg [2:0] state; // @[IFU.scala 55:22]
  reg [127:0] inst_buff; // @[IFU.scala 57:26]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = ~io_reflush_bus_is_reflush; // @[IFU.scala 72:20]
  wire  _T_3 = ~reset; // @[IFU.scala 76:20]
  wire [2:0] _GEN_4 = ~reset ? 3'h1 : state; // @[IFU.scala 76:35 IFU.scala 77:15 IFU.scala 55:22]
  wire [31:0] _GEN_6 = ~reset ? io_reflush_bus_br_target : pc; // @[IFU.scala 76:35 IFU.scala 79:22 IFU.scala 48:16]
  wire  _GEN_8 = ~io_reflush_bus_is_reflush | _T_3; // @[IFU.scala 72:33 IFU.scala 74:23]
  wire [31:0] _GEN_9 = ~io_reflush_bus_is_reflush ? pc : _GEN_6; // @[IFU.scala 72:33 IFU.scala 75:22]
  wire  _GEN_11 = fence_i ? 1'h0 : _GEN_8; // @[IFU.scala 69:20 IFU.scala 71:23]
  wire [31:0] _GEN_12 = fence_i ? pc : _GEN_9; // @[IFU.scala 69:20 IFU.scala 48:16]
  wire  _T_4 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_13 = io_imem_data_ok & ~io_out_ready ? 3'h3 : state; // @[IFU.scala 97:54 IFU.scala 98:15 IFU.scala 55:22]
  wire  _GEN_14 = io_imem_data_ok & ~io_out_ready ? 1'h0 : 1'h1; // @[IFU.scala 97:54 IFU.scala 99:23 IFU.scala 83:21]
  wire [2:0] _GEN_15 = io_imem_data_ok & io_out_ready ? 3'h1 : _GEN_13; // @[IFU.scala 93:53 IFU.scala 94:15]
  wire  _GEN_16 = io_imem_data_ok & io_out_ready | _GEN_14; // @[IFU.scala 93:53 IFU.scala 95:23]
  wire [31:0] _GEN_17 = io_imem_data_ok & io_out_ready ? bp_pc : pc; // @[IFU.scala 93:53 IFU.scala 96:22 IFU.scala 48:16]
  wire [2:0] _GEN_18 = io_reflush_bus_is_reflush & io_imem_data_ok ? 3'h1 : _GEN_15; // @[IFU.scala 89:51 IFU.scala 90:15]
  wire  _GEN_19 = io_reflush_bus_is_reflush & io_imem_data_ok | _GEN_16; // @[IFU.scala 89:51 IFU.scala 91:23]
  wire [31:0] _GEN_20 = io_reflush_bus_is_reflush & io_imem_data_ok ? io_reflush_bus_br_target : _GEN_17; // @[IFU.scala 89:51 IFU.scala 92:22]
  wire [2:0] _GEN_21 = io_reflush_bus_is_reflush & ~io_imem_data_ok ? 3'h2 : _GEN_18; // @[IFU.scala 87:52 IFU.scala 88:15]
  wire  _GEN_22 = io_reflush_bus_is_reflush & ~io_imem_data_ok | _GEN_19; // @[IFU.scala 87:52 IFU.scala 83:21]
  wire [31:0] _GEN_23 = io_reflush_bus_is_reflush & ~io_imem_data_ok ? pc : _GEN_20; // @[IFU.scala 87:52 IFU.scala 48:16]
  wire  _GEN_25 = fence_i ? 1'h0 : _GEN_22; // @[IFU.scala 84:20 IFU.scala 86:23]
  wire [31:0] _GEN_26 = fence_i ? pc : _GEN_23; // @[IFU.scala 84:20 IFU.scala 48:16]
  wire  _T_11 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_27 = io_imem_data_ok ? 3'h1 : state; // @[IFU.scala 106:36 IFU.scala 107:15 IFU.scala 55:22]
  wire [2:0] _GEN_30 = fence_i ? 3'h4 : _GEN_27; // @[IFU.scala 103:20 IFU.scala 104:15]
  wire  _GEN_31 = fence_i ? 1'h0 : io_imem_data_ok; // @[IFU.scala 103:20 IFU.scala 105:23]
  wire  _T_12 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_33 = io_out_ready ? 3'h1 : state; // @[IFU.scala 120:34 IFU.scala 121:15 IFU.scala 55:22]
  wire [31:0] _GEN_35 = io_out_ready ? bp_pc : pc; // @[IFU.scala 120:34 IFU.scala 123:22 IFU.scala 48:16]
  wire [2:0] _GEN_36 = io_reflush_bus_is_reflush ? 3'h1 : _GEN_33; // @[IFU.scala 116:32 IFU.scala 117:15]
  wire  _GEN_37 = io_reflush_bus_is_reflush | io_out_ready; // @[IFU.scala 116:32 IFU.scala 118:23]
  wire [31:0] _GEN_38 = io_reflush_bus_is_reflush ? io_reflush_bus_br_target : _GEN_35; // @[IFU.scala 116:32 IFU.scala 119:22]
  wire [2:0] _GEN_39 = fence_i ? 3'h4 : _GEN_36; // @[IFU.scala 113:20 IFU.scala 114:15]
  wire  _GEN_40 = fence_i ? 1'h0 : _GEN_37; // @[IFU.scala 113:20 IFU.scala 115:23]
  wire [31:0] _GEN_41 = fence_i ? pc : _GEN_38; // @[IFU.scala 113:20 IFU.scala 48:16]
  wire  _T_13 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  icache_fence_finish = io_imem_fence_finish; // @[IFU.scala 33:33 IFU.scala 34:23]
  wire [2:0] _GEN_42 = dcache_fence_finish_0 ? 3'h6 : state; // @[IFU.scala 134:41 IFU.scala 135:15 IFU.scala 55:22]
  wire  _GEN_43 = icache_fence_finish ? 1'h0 : 1'h1; // @[IFU.scala 131:41 IFU.scala 132:23 IFU.scala 127:21]
  wire [2:0] _GEN_44 = icache_fence_finish ? 3'h5 : _GEN_42; // @[IFU.scala 131:41 IFU.scala 133:15]
  wire  _GEN_45 = icache_fence_finish & dcache_fence_finish_0 ? 1'h0 : _GEN_43; // @[IFU.scala 128:57 IFU.scala 129:23]
  wire [2:0] _GEN_46 = icache_fence_finish & dcache_fence_finish_0 ? 3'h0 : _GEN_44; // @[IFU.scala 128:57 IFU.scala 130:15]
  wire  _T_15 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_47 = dcache_fence_finish_0 ? 3'h0 : state; // @[IFU.scala 139:34 IFU.scala 140:15 IFU.scala 55:22]
  wire  _T_16 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_49 = icache_fence_finish ? 3'h0 : state; // @[IFU.scala 144:34 IFU.scala 146:15 IFU.scala 55:22]
  wire [2:0] _GEN_51 = _T_16 ? _GEN_49 : state; // @[Conditional.scala 39:67 IFU.scala 55:22]
  wire [2:0] _GEN_52 = _T_15 ? _GEN_47 : _GEN_51; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_55 = _T_13 ? _GEN_46 : _GEN_52; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_56 = _T_12 ? _GEN_39 : _GEN_55; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_12 & _GEN_40; // @[Conditional.scala 39:67 IFU.scala 47:17]
  wire [31:0] _GEN_58 = _T_12 ? _GEN_41 : pc; // @[Conditional.scala 39:67 IFU.scala 48:16]
  wire  _GEN_59 = _T_12 ? 1'h0 : _T_13 & _GEN_45; // @[Conditional.scala 39:67 IFU.scala 52:17]
  wire  _GEN_61 = _T_11 ? _GEN_31 : _GEN_57; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_62 = _T_11 ? pc : _GEN_58; // @[Conditional.scala 39:67]
  wire  _GEN_63 = _T_11 ? 1'h0 : _GEN_59; // @[Conditional.scala 39:67 IFU.scala 52:17]
  wire  _GEN_64 = _T_4 ? _GEN_25 : _GEN_61; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_66 = _T_4 ? _GEN_26 : _GEN_62; // @[Conditional.scala 39:67]
  wire  _GEN_67 = _T_4 ? 1'h0 : _GEN_63; // @[Conditional.scala 39:67 IFU.scala 52:17]
  reg [2:0] call_count; // @[IFU.scala 151:27]
  reg [2:0] ret_count; // @[IFU.scala 152:26]
  wire  _T_17 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _call_count_T_1 = bp_type == 2'h0 & bp_taken; // @[IFU.scala 158:56]
  wire [2:0] _GEN_77 = {{2'd0}, _call_count_T_1}; // @[IFU.scala 158:30]
  wire [2:0] _call_count_T_3 = call_count + _GEN_77; // @[IFU.scala 158:30]
  wire  _ret_count_T_1 = bp_type == 2'h1 & bp_taken; // @[IFU.scala 159:53]
  wire [2:0] _GEN_78 = {{2'd0}, _ret_count_T_1}; // @[IFU.scala 159:28]
  wire [2:0] _ret_count_T_3 = ret_count + _GEN_78; // @[IFU.scala 159:28]
  wire  _io_out_bits_inst_T_1 = state == 3'h1 & io_imem_data_ok; // @[IFU.scala 179:47]
  wire  _io_out_bits_inst_T_2 = state == 3'h3; // @[IFU.scala 181:15]
  wire [127:0] _io_out_bits_inst_T_3 = state == 3'h3 ? inst_buff : 128'h0; // @[IFU.scala 181:8]
  assign io_imem_valid = _T ? _GEN_11 : _GEN_64; // @[Conditional.scala 40:58]
  assign io_imem_addr = _T ? _GEN_12 : _GEN_66; // @[Conditional.scala 40:58]
  assign io_imem_fence = _T ? 1'h0 : _GEN_67; // @[Conditional.scala 40:58 IFU.scala 52:17]
  assign io_out_valid = _io_out_bits_inst_T_1 & _T_1 | _io_out_bits_inst_T_2 & _T_1; // @[IFU.scala 188:75]
  assign io_out_bits_pc = pc; // @[IFU.scala 178:18]
  assign io_out_bits_inst = state == 3'h1 & io_imem_data_ok ? io_imem_inst : _io_out_bits_inst_T_3; // @[IFU.scala 179:26]
  assign io_out_bits_uncache = ~pc[31]; // @[IFU.scala 175:30]
  assign io_out_bits_offset = pc[3:2]; // @[IFU.scala 176:31]
  assign io_out_bits_bp_br_offset = io_bpu_bp_ok ? io_bpu_bp_offset : bp_offset_reg; // @[IFU.scala 43:19]
  assign io_out_bits_bp_br_taken = io_bpu_bp_ok ? io_bpu_bp_taken : bp_taken_reg; // @[IFU.scala 40:18]
  assign io_out_bits_bp_br_target = io_bpu_bp_ok ? io_bpu_bp_target : bp_pc_reg; // @[IFU.scala 41:15]
  assign io_out_bits_bp_br_type = io_bpu_bp_ok ? io_bpu_bp_type : bp_type_reg; // @[IFU.scala 42:17]
  assign io_bpu_valid = io_imem_valid & (bpu_reg_pc != io_bpu_pc | ~imem_reg_valid); // @[IFU.scala 165:33]
  assign io_bpu_pc = io_imem_addr; // @[IFU.scala 167:13]
  assign io_bpu_is_reflush = io_reflush_bus_is_reflush; // @[IFU.scala 166:21]
  assign io_bpu_call_count = call_count + _GEN_77; // @[IFU.scala 168:35]
  assign io_bpu_ret_count = ret_count + _GEN_78; // @[IFU.scala 169:33]
  assign icache_fence_finish_0 = icache_fence_finish;
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 14:19]
      pc <= 32'h80000000; // @[IFU.scala 14:19]
    end else if (io_reflush_bus_is_reflush) begin // @[IFU.scala 44:12]
      pc <= io_reflush_bus_br_target;
    end else if (io_out_valid & io_out_ready) begin // @[IFU.scala 45:8]
      if (io_bpu_bp_ok) begin // @[IFU.scala 41:15]
        pc <= io_bpu_bp_target;
      end else begin
        pc <= bp_pc_reg;
      end
    end
    if (reset) begin // @[IFU.scala 16:26]
      bp_pc_reg <= 32'h0; // @[IFU.scala 16:26]
    end else if (io_bpu_bp_ok) begin // @[IFU.scala 41:15]
      bp_pc_reg <= io_bpu_bp_target;
    end
    if (reset) begin // @[IFU.scala 18:29]
      bp_taken_reg <= 1'h0; // @[IFU.scala 18:29]
    end else if (io_bpu_bp_ok) begin // @[IFU.scala 40:18]
      bp_taken_reg <= io_bpu_bp_taken;
    end
    if (reset) begin // @[IFU.scala 20:28]
      bp_type_reg <= 2'h0; // @[IFU.scala 20:28]
    end else if (io_bpu_bp_ok) begin // @[IFU.scala 42:17]
      bp_type_reg <= io_bpu_bp_type;
    end
    if (reset) begin // @[IFU.scala 22:30]
      bp_offset_reg <= 2'h0; // @[IFU.scala 22:30]
    end else if (io_bpu_bp_ok) begin // @[IFU.scala 43:19]
      bp_offset_reg <= io_bpu_bp_offset;
    end
    if (reset) begin // @[IFU.scala 24:27]
      bpu_reg_pc <= 32'h0; // @[IFU.scala 24:27]
    end else begin
      bpu_reg_pc <= io_bpu_pc; // @[IFU.scala 162:14]
    end
    if (reset) begin // @[IFU.scala 25:31]
      imem_reg_valid <= 1'h0; // @[IFU.scala 25:31]
    end else begin
      imem_reg_valid <= io_imem_valid; // @[IFU.scala 163:18]
    end
    if (reset) begin // @[IFU.scala 55:22]
      state <= 3'h0; // @[IFU.scala 55:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (fence_i) begin // @[IFU.scala 69:20]
        state <= 3'h4; // @[IFU.scala 70:15]
      end else if (~io_reflush_bus_is_reflush) begin // @[IFU.scala 72:33]
        state <= 3'h1; // @[IFU.scala 73:15]
      end else begin
        state <= _GEN_4;
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      if (fence_i) begin // @[IFU.scala 84:20]
        state <= 3'h4; // @[IFU.scala 85:15]
      end else begin
        state <= _GEN_21;
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      state <= _GEN_30;
    end else begin
      state <= _GEN_56;
    end
    if (reset) begin // @[IFU.scala 57:26]
      inst_buff <= 128'h0; // @[IFU.scala 57:26]
    end else if (io_imem_data_ok) begin // @[IFU.scala 171:26]
      inst_buff <= io_imem_inst; // @[IFU.scala 172:15]
    end
    if (reset) begin // @[IFU.scala 151:27]
      call_count <= 3'h0; // @[IFU.scala 151:27]
    end else if (io_reflush_bus_is_reflush) begin // @[IFU.scala 154:21]
      call_count <= 3'h0; // @[IFU.scala 155:16]
    end else if (_T_17) begin // @[IFU.scala 157:29]
      call_count <= _call_count_T_3; // @[IFU.scala 158:16]
    end
    if (reset) begin // @[IFU.scala 152:26]
      ret_count <= 3'h0; // @[IFU.scala 152:26]
    end else if (io_reflush_bus_is_reflush) begin // @[IFU.scala 154:21]
      ret_count <= 3'h0; // @[IFU.scala 156:15]
    end else if (_T_17) begin // @[IFU.scala 157:29]
      ret_count <= _ret_count_T_3; // @[IFU.scala 159:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  bp_pc_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bp_taken_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bp_type_reg = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  bp_offset_reg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  bpu_reg_pc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  imem_reg_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[2:0];
  _RAND_8 = {4{`RANDOM}};
  inst_buff = _RAND_8[127:0];
  _RAND_9 = {1{`RANDOM}};
  call_count = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  ret_count = _RAND_10[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IQueue(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [31:0]  io_in_bits_pc,
  input  [127:0] io_in_bits_inst,
  input          io_in_bits_uncache,
  input  [1:0]   io_in_bits_offset,
  input  [1:0]   io_in_bits_bp_br_offset,
  input          io_in_bits_bp_br_taken,
  input  [31:0]  io_in_bits_bp_br_target,
  input  [1:0]   io_in_bits_bp_br_type,
  input          io_out_ready,
  output         io_out_valid,
  output         io_out_bits_0_valid,
  output [31:0]  io_out_bits_0_pc,
  output [31:0]  io_out_bits_0_inst,
  output         io_out_bits_0_bp_br_taken,
  output [31:0]  io_out_bits_0_bp_br_target,
  output [1:0]   io_out_bits_0_bp_br_type,
  output         io_out_bits_1_valid,
  output [31:0]  io_out_bits_1_pc,
  output [31:0]  io_out_bits_1_inst,
  output         io_out_bits_1_bp_br_taken,
  output [31:0]  io_out_bits_1_bp_br_target,
  output [1:0]   io_out_bits_1_bp_br_type,
  input          frontend_reflush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] in_counter; // @[IQueue.scala 22:27]
  reg [3:0] out_counter; // @[IQueue.scala 23:28]
  reg [31:0] inst_queue_0_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_0_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_0_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_0_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_0_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_1_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_1_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_1_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_1_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_1_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_2_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_2_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_2_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_2_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_2_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_3_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_3_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_3_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_3_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_3_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_4_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_4_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_4_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_4_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_4_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_5_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_5_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_5_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_5_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_5_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_6_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_6_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_6_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_6_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_6_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_7_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_7_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_7_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_7_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_7_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_8_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_8_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_8_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_8_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_8_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_9_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_9_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_9_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_9_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_9_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_10_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_10_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_10_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_10_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_10_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_11_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_11_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_11_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_11_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_11_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_12_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_12_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_12_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_12_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_12_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_13_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_13_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_13_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_13_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_13_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_14_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_14_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_14_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_14_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_14_bp_br_type; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_15_pc; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_15_inst; // @[IQueue.scala 24:27]
  reg  inst_queue_15_bp_br_taken; // @[IQueue.scala 24:27]
  reg [31:0] inst_queue_15_bp_br_target; // @[IQueue.scala 24:27]
  reg [1:0] inst_queue_15_bp_br_type; // @[IQueue.scala 24:27]
  reg  valid_0; // @[IQueue.scala 26:22]
  reg  valid_1; // @[IQueue.scala 26:22]
  reg  valid_2; // @[IQueue.scala 26:22]
  reg  valid_3; // @[IQueue.scala 26:22]
  reg  valid_4; // @[IQueue.scala 26:22]
  reg  valid_5; // @[IQueue.scala 26:22]
  reg  valid_6; // @[IQueue.scala 26:22]
  reg  valid_7; // @[IQueue.scala 26:22]
  reg  valid_8; // @[IQueue.scala 26:22]
  reg  valid_9; // @[IQueue.scala 26:22]
  reg  valid_10; // @[IQueue.scala 26:22]
  reg  valid_11; // @[IQueue.scala 26:22]
  reg  valid_12; // @[IQueue.scala 26:22]
  reg  valid_13; // @[IQueue.scala 26:22]
  reg  valid_14; // @[IQueue.scala 26:22]
  reg  valid_15; // @[IQueue.scala 26:22]
  wire  has_bp_taken = io_in_bits_bp_br_taken & io_in_bits_offset <= io_in_bits_bp_br_offset; // @[IQueue.scala 30:42]
  wire [1:0] _count_T_2 = 2'h3 - io_in_bits_offset; // @[IQueue.scala 31:35]
  wire [1:0] _count_T_4 = io_in_bits_bp_br_offset - io_in_bits_offset; // @[IQueue.scala 31:80]
  wire [1:0] count = ~has_bp_taken ? _count_T_2 : _count_T_4; // @[IQueue.scala 31:15]
  wire [31:0] in_inst_0 = io_in_bits_inst[31:0]; // @[IQueue.scala 34:32]
  wire [31:0] in_inst_1 = io_in_bits_inst[63:32]; // @[IQueue.scala 35:32]
  wire [31:0] in_inst_2 = io_in_bits_inst[95:64]; // @[IQueue.scala 36:32]
  wire [31:0] in_inst_3 = io_in_bits_inst[127:96]; // @[IQueue.scala 37:32]
  wire [3:0] _full_T_1 = in_counter + 4'h1; // @[IQueue.scala 39:24]
  wire [3:0] _full_T_4 = in_counter + 4'h2; // @[IQueue.scala 39:64]
  wire [3:0] _full_T_8 = in_counter + 4'h3; // @[IQueue.scala 40:18]
  wire  _full_T_9 = _full_T_8 == out_counter; // @[IQueue.scala 40:25]
  wire  _full_T_10 = _full_T_1 == out_counter | _full_T_4 == out_counter | _full_T_9; // @[IQueue.scala 39:88]
  wire [3:0] _full_T_12 = in_counter + 4'h4; // @[IQueue.scala 40:58]
  wire  full = _full_T_10 | _full_T_12 == out_counter; // @[IQueue.scala 40:42]
  wire  _T = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_80 = 4'h0 == in_counter | valid_0; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_81 = 4'h1 == in_counter | valid_1; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_82 = 4'h2 == in_counter | valid_2; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_83 = 4'h3 == in_counter | valid_3; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_84 = 4'h4 == in_counter | valid_4; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_85 = 4'h5 == in_counter | valid_5; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_86 = 4'h6 == in_counter | valid_6; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_87 = 4'h7 == in_counter | valid_7; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_88 = 4'h8 == in_counter | valid_8; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_89 = 4'h9 == in_counter | valid_9; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_90 = 4'ha == in_counter | valid_10; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_91 = 4'hb == in_counter | valid_11; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_92 = 4'hc == in_counter | valid_12; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_93 = 4'hd == in_counter | valid_13; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_94 = 4'he == in_counter | valid_14; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire  _GEN_95 = 4'hf == in_counter | valid_15; // @[IQueue.scala 49:25 IQueue.scala 49:25 IQueue.scala 26:22]
  wire [4:0] _T_2 = {{1'd0}, in_counter}; // @[IQueue.scala 54:33]
  wire [32:0] _inst_queue_pc_T = {{1'd0}, io_in_bits_pc}; // @[IQueue.scala 54:60]
  wire [31:0] _GEN_96 = 4'h0 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_0_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_97 = 4'h1 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_1_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_98 = 4'h2 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_2_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_99 = 4'h3 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_3_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_100 = 4'h4 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_4_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_101 = 4'h5 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_5_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_102 = 4'h6 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_6_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_103 = 4'h7 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_7_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_104 = 4'h8 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_8_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_105 = 4'h9 == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_9_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_106 = 4'ha == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_10_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_107 = 4'hb == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_11_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_108 = 4'hc == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_12_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_109 = 4'hd == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_13_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_110 = 4'he == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_14_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [31:0] _GEN_111 = 4'hf == _T_2[3:0] ? _inst_queue_pc_T[31:0] : inst_queue_15_pc; // @[IQueue.scala 54:43 IQueue.scala 54:43 IQueue.scala 24:27]
  wire [2:0] _inst_queue_inst_T_1 = {{1'd0}, io_in_bits_offset}; // @[IQueue.scala 55:74]
  wire [31:0] _GEN_129 = 2'h1 == _inst_queue_inst_T_1[1:0] ? in_inst_1 : in_inst_0; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_130 = 2'h2 == _inst_queue_inst_T_1[1:0] ? in_inst_2 : _GEN_129; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_131 = 2'h3 == _inst_queue_inst_T_1[1:0] ? in_inst_3 : _GEN_130; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_112 = 4'h0 == _T_2[3:0] ? _GEN_131 : inst_queue_0_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_113 = 4'h1 == _T_2[3:0] ? _GEN_131 : inst_queue_1_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_114 = 4'h2 == _T_2[3:0] ? _GEN_131 : inst_queue_2_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_115 = 4'h3 == _T_2[3:0] ? _GEN_131 : inst_queue_3_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_116 = 4'h4 == _T_2[3:0] ? _GEN_131 : inst_queue_4_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_117 = 4'h5 == _T_2[3:0] ? _GEN_131 : inst_queue_5_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_118 = 4'h6 == _T_2[3:0] ? _GEN_131 : inst_queue_6_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_119 = 4'h7 == _T_2[3:0] ? _GEN_131 : inst_queue_7_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_120 = 4'h8 == _T_2[3:0] ? _GEN_131 : inst_queue_8_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_121 = 4'h9 == _T_2[3:0] ? _GEN_131 : inst_queue_9_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_122 = 4'ha == _T_2[3:0] ? _GEN_131 : inst_queue_10_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_123 = 4'hb == _T_2[3:0] ? _GEN_131 : inst_queue_11_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_124 = 4'hc == _T_2[3:0] ? _GEN_131 : inst_queue_12_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_125 = 4'hd == _T_2[3:0] ? _GEN_131 : inst_queue_13_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_126 = 4'he == _T_2[3:0] ? _GEN_131 : inst_queue_14_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire [31:0] _GEN_127 = 4'hf == _T_2[3:0] ? _GEN_131 : inst_queue_15_inst; // @[IQueue.scala 55:45 IQueue.scala 55:45 IQueue.scala 24:27]
  wire  _GEN_132 = 4'h0 == _T_2[3:0] ? 1'h0 : inst_queue_0_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_133 = 4'h1 == _T_2[3:0] ? 1'h0 : inst_queue_1_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_134 = 4'h2 == _T_2[3:0] ? 1'h0 : inst_queue_2_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_135 = 4'h3 == _T_2[3:0] ? 1'h0 : inst_queue_3_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_136 = 4'h4 == _T_2[3:0] ? 1'h0 : inst_queue_4_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_137 = 4'h5 == _T_2[3:0] ? 1'h0 : inst_queue_5_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_138 = 4'h6 == _T_2[3:0] ? 1'h0 : inst_queue_6_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_139 = 4'h7 == _T_2[3:0] ? 1'h0 : inst_queue_7_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_140 = 4'h8 == _T_2[3:0] ? 1'h0 : inst_queue_8_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_141 = 4'h9 == _T_2[3:0] ? 1'h0 : inst_queue_9_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_142 = 4'ha == _T_2[3:0] ? 1'h0 : inst_queue_10_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_143 = 4'hb == _T_2[3:0] ? 1'h0 : inst_queue_11_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_144 = 4'hc == _T_2[3:0] ? 1'h0 : inst_queue_12_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_145 = 4'hd == _T_2[3:0] ? 1'h0 : inst_queue_13_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_146 = 4'he == _T_2[3:0] ? 1'h0 : inst_queue_14_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire  _GEN_147 = 4'hf == _T_2[3:0] ? 1'h0 : inst_queue_15_bp_br_taken; // @[IQueue.scala 56:52 IQueue.scala 56:52 IQueue.scala 24:27]
  wire [31:0] _GEN_148 = 4'h0 == _T_2[3:0] ? 32'h0 : inst_queue_0_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_149 = 4'h1 == _T_2[3:0] ? 32'h0 : inst_queue_1_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_150 = 4'h2 == _T_2[3:0] ? 32'h0 : inst_queue_2_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_151 = 4'h3 == _T_2[3:0] ? 32'h0 : inst_queue_3_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_152 = 4'h4 == _T_2[3:0] ? 32'h0 : inst_queue_4_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_153 = 4'h5 == _T_2[3:0] ? 32'h0 : inst_queue_5_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_154 = 4'h6 == _T_2[3:0] ? 32'h0 : inst_queue_6_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_155 = 4'h7 == _T_2[3:0] ? 32'h0 : inst_queue_7_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_156 = 4'h8 == _T_2[3:0] ? 32'h0 : inst_queue_8_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_157 = 4'h9 == _T_2[3:0] ? 32'h0 : inst_queue_9_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_158 = 4'ha == _T_2[3:0] ? 32'h0 : inst_queue_10_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_159 = 4'hb == _T_2[3:0] ? 32'h0 : inst_queue_11_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_160 = 4'hc == _T_2[3:0] ? 32'h0 : inst_queue_12_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_161 = 4'hd == _T_2[3:0] ? 32'h0 : inst_queue_13_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_162 = 4'he == _T_2[3:0] ? 32'h0 : inst_queue_14_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [31:0] _GEN_163 = 4'hf == _T_2[3:0] ? 32'h0 : inst_queue_15_bp_br_target; // @[IQueue.scala 57:53 IQueue.scala 57:53 IQueue.scala 24:27]
  wire [1:0] _GEN_164 = 4'h0 == _T_2[3:0] ? 2'h0 : inst_queue_0_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_165 = 4'h1 == _T_2[3:0] ? 2'h0 : inst_queue_1_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_166 = 4'h2 == _T_2[3:0] ? 2'h0 : inst_queue_2_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_167 = 4'h3 == _T_2[3:0] ? 2'h0 : inst_queue_3_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_168 = 4'h4 == _T_2[3:0] ? 2'h0 : inst_queue_4_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_169 = 4'h5 == _T_2[3:0] ? 2'h0 : inst_queue_5_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_170 = 4'h6 == _T_2[3:0] ? 2'h0 : inst_queue_6_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_171 = 4'h7 == _T_2[3:0] ? 2'h0 : inst_queue_7_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_172 = 4'h8 == _T_2[3:0] ? 2'h0 : inst_queue_8_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_173 = 4'h9 == _T_2[3:0] ? 2'h0 : inst_queue_9_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_174 = 4'ha == _T_2[3:0] ? 2'h0 : inst_queue_10_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_175 = 4'hb == _T_2[3:0] ? 2'h0 : inst_queue_11_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_176 = 4'hc == _T_2[3:0] ? 2'h0 : inst_queue_12_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_177 = 4'hd == _T_2[3:0] ? 2'h0 : inst_queue_13_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_178 = 4'he == _T_2[3:0] ? 2'h0 : inst_queue_14_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire [1:0] _GEN_179 = 4'hf == _T_2[3:0] ? 2'h0 : inst_queue_15_bp_br_type; // @[IQueue.scala 58:51 IQueue.scala 58:51 IQueue.scala 24:27]
  wire  _GEN_180 = 4'h0 == _T_2[3:0] | valid_0; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_181 = 4'h1 == _T_2[3:0] | valid_1; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_182 = 4'h2 == _T_2[3:0] | valid_2; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_183 = 4'h3 == _T_2[3:0] | valid_3; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_184 = 4'h4 == _T_2[3:0] | valid_4; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_185 = 4'h5 == _T_2[3:0] | valid_5; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_186 = 4'h6 == _T_2[3:0] | valid_6; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_187 = 4'h7 == _T_2[3:0] | valid_7; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_188 = 4'h8 == _T_2[3:0] | valid_8; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_189 = 4'h9 == _T_2[3:0] | valid_9; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_190 = 4'ha == _T_2[3:0] | valid_10; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_191 = 4'hb == _T_2[3:0] | valid_11; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_192 = 4'hc == _T_2[3:0] | valid_12; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_193 = 4'hd == _T_2[3:0] | valid_13; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_194 = 4'he == _T_2[3:0] | valid_14; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire  _GEN_195 = 4'hf == _T_2[3:0] | valid_15; // @[IQueue.scala 59:35 IQueue.scala 59:35 IQueue.scala 26:22]
  wire [3:0] _GEN_1782 = {{2'd0}, count}; // @[IQueue.scala 62:33]
  wire [3:0] _T_15 = in_counter + _GEN_1782; // @[IQueue.scala 62:33]
  wire  _GEN_292 = 4'h0 == _T_15 ? io_in_bits_bp_br_taken : _GEN_132; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_293 = 4'h1 == _T_15 ? io_in_bits_bp_br_taken : _GEN_133; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_294 = 4'h2 == _T_15 ? io_in_bits_bp_br_taken : _GEN_134; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_295 = 4'h3 == _T_15 ? io_in_bits_bp_br_taken : _GEN_135; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_296 = 4'h4 == _T_15 ? io_in_bits_bp_br_taken : _GEN_136; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_297 = 4'h5 == _T_15 ? io_in_bits_bp_br_taken : _GEN_137; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_298 = 4'h6 == _T_15 ? io_in_bits_bp_br_taken : _GEN_138; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_299 = 4'h7 == _T_15 ? io_in_bits_bp_br_taken : _GEN_139; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_300 = 4'h8 == _T_15 ? io_in_bits_bp_br_taken : _GEN_140; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_301 = 4'h9 == _T_15 ? io_in_bits_bp_br_taken : _GEN_141; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_302 = 4'ha == _T_15 ? io_in_bits_bp_br_taken : _GEN_142; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_303 = 4'hb == _T_15 ? io_in_bits_bp_br_taken : _GEN_143; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_304 = 4'hc == _T_15 ? io_in_bits_bp_br_taken : _GEN_144; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_305 = 4'hd == _T_15 ? io_in_bits_bp_br_taken : _GEN_145; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_306 = 4'he == _T_15 ? io_in_bits_bp_br_taken : _GEN_146; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_307 = 4'hf == _T_15 ? io_in_bits_bp_br_taken : _GEN_147; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire [31:0] _GEN_308 = 4'h0 == _T_15 ? io_in_bits_bp_br_target : _GEN_148; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_309 = 4'h1 == _T_15 ? io_in_bits_bp_br_target : _GEN_149; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_310 = 4'h2 == _T_15 ? io_in_bits_bp_br_target : _GEN_150; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_311 = 4'h3 == _T_15 ? io_in_bits_bp_br_target : _GEN_151; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_312 = 4'h4 == _T_15 ? io_in_bits_bp_br_target : _GEN_152; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_313 = 4'h5 == _T_15 ? io_in_bits_bp_br_target : _GEN_153; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_314 = 4'h6 == _T_15 ? io_in_bits_bp_br_target : _GEN_154; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_315 = 4'h7 == _T_15 ? io_in_bits_bp_br_target : _GEN_155; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_316 = 4'h8 == _T_15 ? io_in_bits_bp_br_target : _GEN_156; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_317 = 4'h9 == _T_15 ? io_in_bits_bp_br_target : _GEN_157; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_318 = 4'ha == _T_15 ? io_in_bits_bp_br_target : _GEN_158; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_319 = 4'hb == _T_15 ? io_in_bits_bp_br_target : _GEN_159; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_320 = 4'hc == _T_15 ? io_in_bits_bp_br_target : _GEN_160; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_321 = 4'hd == _T_15 ? io_in_bits_bp_br_target : _GEN_161; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_322 = 4'he == _T_15 ? io_in_bits_bp_br_target : _GEN_162; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_323 = 4'hf == _T_15 ? io_in_bits_bp_br_target : _GEN_163; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [1:0] _GEN_324 = 4'h0 == _T_15 ? io_in_bits_bp_br_type : _GEN_164; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_325 = 4'h1 == _T_15 ? io_in_bits_bp_br_type : _GEN_165; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_326 = 4'h2 == _T_15 ? io_in_bits_bp_br_type : _GEN_166; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_327 = 4'h3 == _T_15 ? io_in_bits_bp_br_type : _GEN_167; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_328 = 4'h4 == _T_15 ? io_in_bits_bp_br_type : _GEN_168; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_329 = 4'h5 == _T_15 ? io_in_bits_bp_br_type : _GEN_169; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_330 = 4'h6 == _T_15 ? io_in_bits_bp_br_type : _GEN_170; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_331 = 4'h7 == _T_15 ? io_in_bits_bp_br_type : _GEN_171; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_332 = 4'h8 == _T_15 ? io_in_bits_bp_br_type : _GEN_172; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_333 = 4'h9 == _T_15 ? io_in_bits_bp_br_type : _GEN_173; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_334 = 4'ha == _T_15 ? io_in_bits_bp_br_type : _GEN_174; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_335 = 4'hb == _T_15 ? io_in_bits_bp_br_type : _GEN_175; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_336 = 4'hc == _T_15 ? io_in_bits_bp_br_type : _GEN_176; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_337 = 4'hd == _T_15 ? io_in_bits_bp_br_type : _GEN_177; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_338 = 4'he == _T_15 ? io_in_bits_bp_br_type : _GEN_178; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_339 = 4'hf == _T_15 ? io_in_bits_bp_br_type : _GEN_179; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire  _GEN_340 = has_bp_taken ? _GEN_292 : _GEN_132; // @[IQueue.scala 61:29]
  wire  _GEN_341 = has_bp_taken ? _GEN_293 : _GEN_133; // @[IQueue.scala 61:29]
  wire  _GEN_342 = has_bp_taken ? _GEN_294 : _GEN_134; // @[IQueue.scala 61:29]
  wire  _GEN_343 = has_bp_taken ? _GEN_295 : _GEN_135; // @[IQueue.scala 61:29]
  wire  _GEN_344 = has_bp_taken ? _GEN_296 : _GEN_136; // @[IQueue.scala 61:29]
  wire  _GEN_345 = has_bp_taken ? _GEN_297 : _GEN_137; // @[IQueue.scala 61:29]
  wire  _GEN_346 = has_bp_taken ? _GEN_298 : _GEN_138; // @[IQueue.scala 61:29]
  wire  _GEN_347 = has_bp_taken ? _GEN_299 : _GEN_139; // @[IQueue.scala 61:29]
  wire  _GEN_348 = has_bp_taken ? _GEN_300 : _GEN_140; // @[IQueue.scala 61:29]
  wire  _GEN_349 = has_bp_taken ? _GEN_301 : _GEN_141; // @[IQueue.scala 61:29]
  wire  _GEN_350 = has_bp_taken ? _GEN_302 : _GEN_142; // @[IQueue.scala 61:29]
  wire  _GEN_351 = has_bp_taken ? _GEN_303 : _GEN_143; // @[IQueue.scala 61:29]
  wire  _GEN_352 = has_bp_taken ? _GEN_304 : _GEN_144; // @[IQueue.scala 61:29]
  wire  _GEN_353 = has_bp_taken ? _GEN_305 : _GEN_145; // @[IQueue.scala 61:29]
  wire  _GEN_354 = has_bp_taken ? _GEN_306 : _GEN_146; // @[IQueue.scala 61:29]
  wire  _GEN_355 = has_bp_taken ? _GEN_307 : _GEN_147; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_356 = has_bp_taken ? _GEN_308 : _GEN_148; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_357 = has_bp_taken ? _GEN_309 : _GEN_149; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_358 = has_bp_taken ? _GEN_310 : _GEN_150; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_359 = has_bp_taken ? _GEN_311 : _GEN_151; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_360 = has_bp_taken ? _GEN_312 : _GEN_152; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_361 = has_bp_taken ? _GEN_313 : _GEN_153; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_362 = has_bp_taken ? _GEN_314 : _GEN_154; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_363 = has_bp_taken ? _GEN_315 : _GEN_155; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_364 = has_bp_taken ? _GEN_316 : _GEN_156; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_365 = has_bp_taken ? _GEN_317 : _GEN_157; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_366 = has_bp_taken ? _GEN_318 : _GEN_158; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_367 = has_bp_taken ? _GEN_319 : _GEN_159; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_368 = has_bp_taken ? _GEN_320 : _GEN_160; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_369 = has_bp_taken ? _GEN_321 : _GEN_161; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_370 = has_bp_taken ? _GEN_322 : _GEN_162; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_371 = has_bp_taken ? _GEN_323 : _GEN_163; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_372 = has_bp_taken ? _GEN_324 : _GEN_164; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_373 = has_bp_taken ? _GEN_325 : _GEN_165; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_374 = has_bp_taken ? _GEN_326 : _GEN_166; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_375 = has_bp_taken ? _GEN_327 : _GEN_167; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_376 = has_bp_taken ? _GEN_328 : _GEN_168; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_377 = has_bp_taken ? _GEN_329 : _GEN_169; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_378 = has_bp_taken ? _GEN_330 : _GEN_170; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_379 = has_bp_taken ? _GEN_331 : _GEN_171; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_380 = has_bp_taken ? _GEN_332 : _GEN_172; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_381 = has_bp_taken ? _GEN_333 : _GEN_173; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_382 = has_bp_taken ? _GEN_334 : _GEN_174; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_383 = has_bp_taken ? _GEN_335 : _GEN_175; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_384 = has_bp_taken ? _GEN_336 : _GEN_176; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_385 = has_bp_taken ? _GEN_337 : _GEN_177; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_386 = has_bp_taken ? _GEN_338 : _GEN_178; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_387 = has_bp_taken ? _GEN_339 : _GEN_179; // @[IQueue.scala 61:29]
  wire [3:0] _in_counter_T_5 = _T_15 + 4'h1; // @[IQueue.scala 66:44]
  wire [31:0] _inst_queue_pc_T_3 = io_in_bits_pc + 32'h4; // @[IQueue.scala 54:60]
  wire [31:0] _GEN_388 = 4'h0 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_96; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_389 = 4'h1 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_97; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_390 = 4'h2 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_98; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_391 = 4'h3 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_99; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_392 = 4'h4 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_100; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_393 = 4'h5 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_101; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_394 = 4'h6 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_102; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_395 = 4'h7 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_103; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_396 = 4'h8 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_104; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_397 = 4'h9 == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_105; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_398 = 4'ha == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_106; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_399 = 4'hb == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_107; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_400 = 4'hc == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_108; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_401 = 4'hd == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_109; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_402 = 4'he == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_110; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_403 = 4'hf == _full_T_1 ? _inst_queue_pc_T_3 : _GEN_111; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [1:0] _inst_queue_inst_T_4 = io_in_bits_offset + 2'h1; // @[IQueue.scala 55:74]
  wire [31:0] _GEN_421 = 2'h1 == _inst_queue_inst_T_4 ? in_inst_1 : in_inst_0; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_422 = 2'h2 == _inst_queue_inst_T_4 ? in_inst_2 : _GEN_421; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_423 = 2'h3 == _inst_queue_inst_T_4 ? in_inst_3 : _GEN_422; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_404 = 4'h0 == _full_T_1 ? _GEN_423 : _GEN_112; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_405 = 4'h1 == _full_T_1 ? _GEN_423 : _GEN_113; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_406 = 4'h2 == _full_T_1 ? _GEN_423 : _GEN_114; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_407 = 4'h3 == _full_T_1 ? _GEN_423 : _GEN_115; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_408 = 4'h4 == _full_T_1 ? _GEN_423 : _GEN_116; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_409 = 4'h5 == _full_T_1 ? _GEN_423 : _GEN_117; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_410 = 4'h6 == _full_T_1 ? _GEN_423 : _GEN_118; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_411 = 4'h7 == _full_T_1 ? _GEN_423 : _GEN_119; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_412 = 4'h8 == _full_T_1 ? _GEN_423 : _GEN_120; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_413 = 4'h9 == _full_T_1 ? _GEN_423 : _GEN_121; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_414 = 4'ha == _full_T_1 ? _GEN_423 : _GEN_122; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_415 = 4'hb == _full_T_1 ? _GEN_423 : _GEN_123; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_416 = 4'hc == _full_T_1 ? _GEN_423 : _GEN_124; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_417 = 4'hd == _full_T_1 ? _GEN_423 : _GEN_125; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_418 = 4'he == _full_T_1 ? _GEN_423 : _GEN_126; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_419 = 4'hf == _full_T_1 ? _GEN_423 : _GEN_127; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire  _GEN_424 = 4'h0 == _full_T_1 ? 1'h0 : _GEN_340; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_425 = 4'h1 == _full_T_1 ? 1'h0 : _GEN_341; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_426 = 4'h2 == _full_T_1 ? 1'h0 : _GEN_342; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_427 = 4'h3 == _full_T_1 ? 1'h0 : _GEN_343; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_428 = 4'h4 == _full_T_1 ? 1'h0 : _GEN_344; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_429 = 4'h5 == _full_T_1 ? 1'h0 : _GEN_345; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_430 = 4'h6 == _full_T_1 ? 1'h0 : _GEN_346; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_431 = 4'h7 == _full_T_1 ? 1'h0 : _GEN_347; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_432 = 4'h8 == _full_T_1 ? 1'h0 : _GEN_348; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_433 = 4'h9 == _full_T_1 ? 1'h0 : _GEN_349; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_434 = 4'ha == _full_T_1 ? 1'h0 : _GEN_350; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_435 = 4'hb == _full_T_1 ? 1'h0 : _GEN_351; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_436 = 4'hc == _full_T_1 ? 1'h0 : _GEN_352; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_437 = 4'hd == _full_T_1 ? 1'h0 : _GEN_353; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_438 = 4'he == _full_T_1 ? 1'h0 : _GEN_354; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_439 = 4'hf == _full_T_1 ? 1'h0 : _GEN_355; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire [31:0] _GEN_440 = 4'h0 == _full_T_1 ? 32'h0 : _GEN_356; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_441 = 4'h1 == _full_T_1 ? 32'h0 : _GEN_357; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_442 = 4'h2 == _full_T_1 ? 32'h0 : _GEN_358; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_443 = 4'h3 == _full_T_1 ? 32'h0 : _GEN_359; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_444 = 4'h4 == _full_T_1 ? 32'h0 : _GEN_360; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_445 = 4'h5 == _full_T_1 ? 32'h0 : _GEN_361; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_446 = 4'h6 == _full_T_1 ? 32'h0 : _GEN_362; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_447 = 4'h7 == _full_T_1 ? 32'h0 : _GEN_363; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_448 = 4'h8 == _full_T_1 ? 32'h0 : _GEN_364; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_449 = 4'h9 == _full_T_1 ? 32'h0 : _GEN_365; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_450 = 4'ha == _full_T_1 ? 32'h0 : _GEN_366; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_451 = 4'hb == _full_T_1 ? 32'h0 : _GEN_367; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_452 = 4'hc == _full_T_1 ? 32'h0 : _GEN_368; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_453 = 4'hd == _full_T_1 ? 32'h0 : _GEN_369; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_454 = 4'he == _full_T_1 ? 32'h0 : _GEN_370; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_455 = 4'hf == _full_T_1 ? 32'h0 : _GEN_371; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [1:0] _GEN_456 = 4'h0 == _full_T_1 ? 2'h0 : _GEN_372; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_457 = 4'h1 == _full_T_1 ? 2'h0 : _GEN_373; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_458 = 4'h2 == _full_T_1 ? 2'h0 : _GEN_374; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_459 = 4'h3 == _full_T_1 ? 2'h0 : _GEN_375; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_460 = 4'h4 == _full_T_1 ? 2'h0 : _GEN_376; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_461 = 4'h5 == _full_T_1 ? 2'h0 : _GEN_377; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_462 = 4'h6 == _full_T_1 ? 2'h0 : _GEN_378; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_463 = 4'h7 == _full_T_1 ? 2'h0 : _GEN_379; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_464 = 4'h8 == _full_T_1 ? 2'h0 : _GEN_380; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_465 = 4'h9 == _full_T_1 ? 2'h0 : _GEN_381; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_466 = 4'ha == _full_T_1 ? 2'h0 : _GEN_382; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_467 = 4'hb == _full_T_1 ? 2'h0 : _GEN_383; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_468 = 4'hc == _full_T_1 ? 2'h0 : _GEN_384; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_469 = 4'hd == _full_T_1 ? 2'h0 : _GEN_385; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_470 = 4'he == _full_T_1 ? 2'h0 : _GEN_386; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_471 = 4'hf == _full_T_1 ? 2'h0 : _GEN_387; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire  _GEN_472 = 4'h0 == _full_T_1 | _GEN_180; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_473 = 4'h1 == _full_T_1 | _GEN_181; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_474 = 4'h2 == _full_T_1 | _GEN_182; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_475 = 4'h3 == _full_T_1 | _GEN_183; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_476 = 4'h4 == _full_T_1 | _GEN_184; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_477 = 4'h5 == _full_T_1 | _GEN_185; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_478 = 4'h6 == _full_T_1 | _GEN_186; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_479 = 4'h7 == _full_T_1 | _GEN_187; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_480 = 4'h8 == _full_T_1 | _GEN_188; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_481 = 4'h9 == _full_T_1 | _GEN_189; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_482 = 4'ha == _full_T_1 | _GEN_190; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_483 = 4'hb == _full_T_1 | _GEN_191; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_484 = 4'hc == _full_T_1 | _GEN_192; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_485 = 4'hd == _full_T_1 | _GEN_193; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_486 = 4'he == _full_T_1 | _GEN_194; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_487 = 4'hf == _full_T_1 | _GEN_195; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire [31:0] _GEN_488 = 2'h1 <= count ? _GEN_388 : _GEN_96; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_489 = 2'h1 <= count ? _GEN_389 : _GEN_97; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_490 = 2'h1 <= count ? _GEN_390 : _GEN_98; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_491 = 2'h1 <= count ? _GEN_391 : _GEN_99; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_492 = 2'h1 <= count ? _GEN_392 : _GEN_100; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_493 = 2'h1 <= count ? _GEN_393 : _GEN_101; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_494 = 2'h1 <= count ? _GEN_394 : _GEN_102; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_495 = 2'h1 <= count ? _GEN_395 : _GEN_103; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_496 = 2'h1 <= count ? _GEN_396 : _GEN_104; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_497 = 2'h1 <= count ? _GEN_397 : _GEN_105; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_498 = 2'h1 <= count ? _GEN_398 : _GEN_106; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_499 = 2'h1 <= count ? _GEN_399 : _GEN_107; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_500 = 2'h1 <= count ? _GEN_400 : _GEN_108; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_501 = 2'h1 <= count ? _GEN_401 : _GEN_109; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_502 = 2'h1 <= count ? _GEN_402 : _GEN_110; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_503 = 2'h1 <= count ? _GEN_403 : _GEN_111; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_504 = 2'h1 <= count ? _GEN_404 : _GEN_112; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_505 = 2'h1 <= count ? _GEN_405 : _GEN_113; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_506 = 2'h1 <= count ? _GEN_406 : _GEN_114; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_507 = 2'h1 <= count ? _GEN_407 : _GEN_115; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_508 = 2'h1 <= count ? _GEN_408 : _GEN_116; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_509 = 2'h1 <= count ? _GEN_409 : _GEN_117; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_510 = 2'h1 <= count ? _GEN_410 : _GEN_118; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_511 = 2'h1 <= count ? _GEN_411 : _GEN_119; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_512 = 2'h1 <= count ? _GEN_412 : _GEN_120; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_513 = 2'h1 <= count ? _GEN_413 : _GEN_121; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_514 = 2'h1 <= count ? _GEN_414 : _GEN_122; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_515 = 2'h1 <= count ? _GEN_415 : _GEN_123; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_516 = 2'h1 <= count ? _GEN_416 : _GEN_124; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_517 = 2'h1 <= count ? _GEN_417 : _GEN_125; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_518 = 2'h1 <= count ? _GEN_418 : _GEN_126; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_519 = 2'h1 <= count ? _GEN_419 : _GEN_127; // @[IQueue.scala 53:29]
  wire  _GEN_520 = 2'h1 <= count ? _GEN_424 : _GEN_340; // @[IQueue.scala 53:29]
  wire  _GEN_521 = 2'h1 <= count ? _GEN_425 : _GEN_341; // @[IQueue.scala 53:29]
  wire  _GEN_522 = 2'h1 <= count ? _GEN_426 : _GEN_342; // @[IQueue.scala 53:29]
  wire  _GEN_523 = 2'h1 <= count ? _GEN_427 : _GEN_343; // @[IQueue.scala 53:29]
  wire  _GEN_524 = 2'h1 <= count ? _GEN_428 : _GEN_344; // @[IQueue.scala 53:29]
  wire  _GEN_525 = 2'h1 <= count ? _GEN_429 : _GEN_345; // @[IQueue.scala 53:29]
  wire  _GEN_526 = 2'h1 <= count ? _GEN_430 : _GEN_346; // @[IQueue.scala 53:29]
  wire  _GEN_527 = 2'h1 <= count ? _GEN_431 : _GEN_347; // @[IQueue.scala 53:29]
  wire  _GEN_528 = 2'h1 <= count ? _GEN_432 : _GEN_348; // @[IQueue.scala 53:29]
  wire  _GEN_529 = 2'h1 <= count ? _GEN_433 : _GEN_349; // @[IQueue.scala 53:29]
  wire  _GEN_530 = 2'h1 <= count ? _GEN_434 : _GEN_350; // @[IQueue.scala 53:29]
  wire  _GEN_531 = 2'h1 <= count ? _GEN_435 : _GEN_351; // @[IQueue.scala 53:29]
  wire  _GEN_532 = 2'h1 <= count ? _GEN_436 : _GEN_352; // @[IQueue.scala 53:29]
  wire  _GEN_533 = 2'h1 <= count ? _GEN_437 : _GEN_353; // @[IQueue.scala 53:29]
  wire  _GEN_534 = 2'h1 <= count ? _GEN_438 : _GEN_354; // @[IQueue.scala 53:29]
  wire  _GEN_535 = 2'h1 <= count ? _GEN_439 : _GEN_355; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_536 = 2'h1 <= count ? _GEN_440 : _GEN_356; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_537 = 2'h1 <= count ? _GEN_441 : _GEN_357; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_538 = 2'h1 <= count ? _GEN_442 : _GEN_358; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_539 = 2'h1 <= count ? _GEN_443 : _GEN_359; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_540 = 2'h1 <= count ? _GEN_444 : _GEN_360; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_541 = 2'h1 <= count ? _GEN_445 : _GEN_361; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_542 = 2'h1 <= count ? _GEN_446 : _GEN_362; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_543 = 2'h1 <= count ? _GEN_447 : _GEN_363; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_544 = 2'h1 <= count ? _GEN_448 : _GEN_364; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_545 = 2'h1 <= count ? _GEN_449 : _GEN_365; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_546 = 2'h1 <= count ? _GEN_450 : _GEN_366; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_547 = 2'h1 <= count ? _GEN_451 : _GEN_367; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_548 = 2'h1 <= count ? _GEN_452 : _GEN_368; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_549 = 2'h1 <= count ? _GEN_453 : _GEN_369; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_550 = 2'h1 <= count ? _GEN_454 : _GEN_370; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_551 = 2'h1 <= count ? _GEN_455 : _GEN_371; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_552 = 2'h1 <= count ? _GEN_456 : _GEN_372; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_553 = 2'h1 <= count ? _GEN_457 : _GEN_373; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_554 = 2'h1 <= count ? _GEN_458 : _GEN_374; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_555 = 2'h1 <= count ? _GEN_459 : _GEN_375; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_556 = 2'h1 <= count ? _GEN_460 : _GEN_376; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_557 = 2'h1 <= count ? _GEN_461 : _GEN_377; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_558 = 2'h1 <= count ? _GEN_462 : _GEN_378; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_559 = 2'h1 <= count ? _GEN_463 : _GEN_379; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_560 = 2'h1 <= count ? _GEN_464 : _GEN_380; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_561 = 2'h1 <= count ? _GEN_465 : _GEN_381; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_562 = 2'h1 <= count ? _GEN_466 : _GEN_382; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_563 = 2'h1 <= count ? _GEN_467 : _GEN_383; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_564 = 2'h1 <= count ? _GEN_468 : _GEN_384; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_565 = 2'h1 <= count ? _GEN_469 : _GEN_385; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_566 = 2'h1 <= count ? _GEN_470 : _GEN_386; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_567 = 2'h1 <= count ? _GEN_471 : _GEN_387; // @[IQueue.scala 53:29]
  wire  _GEN_568 = 2'h1 <= count ? _GEN_472 : _GEN_180; // @[IQueue.scala 53:29]
  wire  _GEN_569 = 2'h1 <= count ? _GEN_473 : _GEN_181; // @[IQueue.scala 53:29]
  wire  _GEN_570 = 2'h1 <= count ? _GEN_474 : _GEN_182; // @[IQueue.scala 53:29]
  wire  _GEN_571 = 2'h1 <= count ? _GEN_475 : _GEN_183; // @[IQueue.scala 53:29]
  wire  _GEN_572 = 2'h1 <= count ? _GEN_476 : _GEN_184; // @[IQueue.scala 53:29]
  wire  _GEN_573 = 2'h1 <= count ? _GEN_477 : _GEN_185; // @[IQueue.scala 53:29]
  wire  _GEN_574 = 2'h1 <= count ? _GEN_478 : _GEN_186; // @[IQueue.scala 53:29]
  wire  _GEN_575 = 2'h1 <= count ? _GEN_479 : _GEN_187; // @[IQueue.scala 53:29]
  wire  _GEN_576 = 2'h1 <= count ? _GEN_480 : _GEN_188; // @[IQueue.scala 53:29]
  wire  _GEN_577 = 2'h1 <= count ? _GEN_481 : _GEN_189; // @[IQueue.scala 53:29]
  wire  _GEN_578 = 2'h1 <= count ? _GEN_482 : _GEN_190; // @[IQueue.scala 53:29]
  wire  _GEN_579 = 2'h1 <= count ? _GEN_483 : _GEN_191; // @[IQueue.scala 53:29]
  wire  _GEN_580 = 2'h1 <= count ? _GEN_484 : _GEN_192; // @[IQueue.scala 53:29]
  wire  _GEN_581 = 2'h1 <= count ? _GEN_485 : _GEN_193; // @[IQueue.scala 53:29]
  wire  _GEN_582 = 2'h1 <= count ? _GEN_486 : _GEN_194; // @[IQueue.scala 53:29]
  wire  _GEN_583 = 2'h1 <= count ? _GEN_487 : _GEN_195; // @[IQueue.scala 53:29]
  wire  _GEN_584 = 4'h0 == _T_15 ? io_in_bits_bp_br_taken : _GEN_520; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_585 = 4'h1 == _T_15 ? io_in_bits_bp_br_taken : _GEN_521; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_586 = 4'h2 == _T_15 ? io_in_bits_bp_br_taken : _GEN_522; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_587 = 4'h3 == _T_15 ? io_in_bits_bp_br_taken : _GEN_523; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_588 = 4'h4 == _T_15 ? io_in_bits_bp_br_taken : _GEN_524; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_589 = 4'h5 == _T_15 ? io_in_bits_bp_br_taken : _GEN_525; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_590 = 4'h6 == _T_15 ? io_in_bits_bp_br_taken : _GEN_526; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_591 = 4'h7 == _T_15 ? io_in_bits_bp_br_taken : _GEN_527; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_592 = 4'h8 == _T_15 ? io_in_bits_bp_br_taken : _GEN_528; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_593 = 4'h9 == _T_15 ? io_in_bits_bp_br_taken : _GEN_529; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_594 = 4'ha == _T_15 ? io_in_bits_bp_br_taken : _GEN_530; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_595 = 4'hb == _T_15 ? io_in_bits_bp_br_taken : _GEN_531; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_596 = 4'hc == _T_15 ? io_in_bits_bp_br_taken : _GEN_532; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_597 = 4'hd == _T_15 ? io_in_bits_bp_br_taken : _GEN_533; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_598 = 4'he == _T_15 ? io_in_bits_bp_br_taken : _GEN_534; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_599 = 4'hf == _T_15 ? io_in_bits_bp_br_taken : _GEN_535; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire [31:0] _GEN_600 = 4'h0 == _T_15 ? io_in_bits_bp_br_target : _GEN_536; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_601 = 4'h1 == _T_15 ? io_in_bits_bp_br_target : _GEN_537; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_602 = 4'h2 == _T_15 ? io_in_bits_bp_br_target : _GEN_538; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_603 = 4'h3 == _T_15 ? io_in_bits_bp_br_target : _GEN_539; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_604 = 4'h4 == _T_15 ? io_in_bits_bp_br_target : _GEN_540; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_605 = 4'h5 == _T_15 ? io_in_bits_bp_br_target : _GEN_541; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_606 = 4'h6 == _T_15 ? io_in_bits_bp_br_target : _GEN_542; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_607 = 4'h7 == _T_15 ? io_in_bits_bp_br_target : _GEN_543; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_608 = 4'h8 == _T_15 ? io_in_bits_bp_br_target : _GEN_544; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_609 = 4'h9 == _T_15 ? io_in_bits_bp_br_target : _GEN_545; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_610 = 4'ha == _T_15 ? io_in_bits_bp_br_target : _GEN_546; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_611 = 4'hb == _T_15 ? io_in_bits_bp_br_target : _GEN_547; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_612 = 4'hc == _T_15 ? io_in_bits_bp_br_target : _GEN_548; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_613 = 4'hd == _T_15 ? io_in_bits_bp_br_target : _GEN_549; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_614 = 4'he == _T_15 ? io_in_bits_bp_br_target : _GEN_550; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_615 = 4'hf == _T_15 ? io_in_bits_bp_br_target : _GEN_551; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [1:0] _GEN_616 = 4'h0 == _T_15 ? io_in_bits_bp_br_type : _GEN_552; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_617 = 4'h1 == _T_15 ? io_in_bits_bp_br_type : _GEN_553; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_618 = 4'h2 == _T_15 ? io_in_bits_bp_br_type : _GEN_554; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_619 = 4'h3 == _T_15 ? io_in_bits_bp_br_type : _GEN_555; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_620 = 4'h4 == _T_15 ? io_in_bits_bp_br_type : _GEN_556; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_621 = 4'h5 == _T_15 ? io_in_bits_bp_br_type : _GEN_557; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_622 = 4'h6 == _T_15 ? io_in_bits_bp_br_type : _GEN_558; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_623 = 4'h7 == _T_15 ? io_in_bits_bp_br_type : _GEN_559; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_624 = 4'h8 == _T_15 ? io_in_bits_bp_br_type : _GEN_560; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_625 = 4'h9 == _T_15 ? io_in_bits_bp_br_type : _GEN_561; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_626 = 4'ha == _T_15 ? io_in_bits_bp_br_type : _GEN_562; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_627 = 4'hb == _T_15 ? io_in_bits_bp_br_type : _GEN_563; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_628 = 4'hc == _T_15 ? io_in_bits_bp_br_type : _GEN_564; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_629 = 4'hd == _T_15 ? io_in_bits_bp_br_type : _GEN_565; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_630 = 4'he == _T_15 ? io_in_bits_bp_br_type : _GEN_566; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_631 = 4'hf == _T_15 ? io_in_bits_bp_br_type : _GEN_567; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire  _GEN_632 = has_bp_taken ? _GEN_584 : _GEN_520; // @[IQueue.scala 61:29]
  wire  _GEN_633 = has_bp_taken ? _GEN_585 : _GEN_521; // @[IQueue.scala 61:29]
  wire  _GEN_634 = has_bp_taken ? _GEN_586 : _GEN_522; // @[IQueue.scala 61:29]
  wire  _GEN_635 = has_bp_taken ? _GEN_587 : _GEN_523; // @[IQueue.scala 61:29]
  wire  _GEN_636 = has_bp_taken ? _GEN_588 : _GEN_524; // @[IQueue.scala 61:29]
  wire  _GEN_637 = has_bp_taken ? _GEN_589 : _GEN_525; // @[IQueue.scala 61:29]
  wire  _GEN_638 = has_bp_taken ? _GEN_590 : _GEN_526; // @[IQueue.scala 61:29]
  wire  _GEN_639 = has_bp_taken ? _GEN_591 : _GEN_527; // @[IQueue.scala 61:29]
  wire  _GEN_640 = has_bp_taken ? _GEN_592 : _GEN_528; // @[IQueue.scala 61:29]
  wire  _GEN_641 = has_bp_taken ? _GEN_593 : _GEN_529; // @[IQueue.scala 61:29]
  wire  _GEN_642 = has_bp_taken ? _GEN_594 : _GEN_530; // @[IQueue.scala 61:29]
  wire  _GEN_643 = has_bp_taken ? _GEN_595 : _GEN_531; // @[IQueue.scala 61:29]
  wire  _GEN_644 = has_bp_taken ? _GEN_596 : _GEN_532; // @[IQueue.scala 61:29]
  wire  _GEN_645 = has_bp_taken ? _GEN_597 : _GEN_533; // @[IQueue.scala 61:29]
  wire  _GEN_646 = has_bp_taken ? _GEN_598 : _GEN_534; // @[IQueue.scala 61:29]
  wire  _GEN_647 = has_bp_taken ? _GEN_599 : _GEN_535; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_648 = has_bp_taken ? _GEN_600 : _GEN_536; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_649 = has_bp_taken ? _GEN_601 : _GEN_537; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_650 = has_bp_taken ? _GEN_602 : _GEN_538; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_651 = has_bp_taken ? _GEN_603 : _GEN_539; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_652 = has_bp_taken ? _GEN_604 : _GEN_540; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_653 = has_bp_taken ? _GEN_605 : _GEN_541; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_654 = has_bp_taken ? _GEN_606 : _GEN_542; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_655 = has_bp_taken ? _GEN_607 : _GEN_543; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_656 = has_bp_taken ? _GEN_608 : _GEN_544; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_657 = has_bp_taken ? _GEN_609 : _GEN_545; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_658 = has_bp_taken ? _GEN_610 : _GEN_546; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_659 = has_bp_taken ? _GEN_611 : _GEN_547; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_660 = has_bp_taken ? _GEN_612 : _GEN_548; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_661 = has_bp_taken ? _GEN_613 : _GEN_549; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_662 = has_bp_taken ? _GEN_614 : _GEN_550; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_663 = has_bp_taken ? _GEN_615 : _GEN_551; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_664 = has_bp_taken ? _GEN_616 : _GEN_552; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_665 = has_bp_taken ? _GEN_617 : _GEN_553; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_666 = has_bp_taken ? _GEN_618 : _GEN_554; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_667 = has_bp_taken ? _GEN_619 : _GEN_555; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_668 = has_bp_taken ? _GEN_620 : _GEN_556; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_669 = has_bp_taken ? _GEN_621 : _GEN_557; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_670 = has_bp_taken ? _GEN_622 : _GEN_558; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_671 = has_bp_taken ? _GEN_623 : _GEN_559; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_672 = has_bp_taken ? _GEN_624 : _GEN_560; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_673 = has_bp_taken ? _GEN_625 : _GEN_561; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_674 = has_bp_taken ? _GEN_626 : _GEN_562; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_675 = has_bp_taken ? _GEN_627 : _GEN_563; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_676 = has_bp_taken ? _GEN_628 : _GEN_564; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_677 = has_bp_taken ? _GEN_629 : _GEN_565; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_678 = has_bp_taken ? _GEN_630 : _GEN_566; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_679 = has_bp_taken ? _GEN_631 : _GEN_567; // @[IQueue.scala 61:29]
  wire [31:0] _inst_queue_pc_T_5 = io_in_bits_pc + 32'h8; // @[IQueue.scala 54:60]
  wire [31:0] _GEN_680 = 4'h0 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_488; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_681 = 4'h1 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_489; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_682 = 4'h2 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_490; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_683 = 4'h3 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_491; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_684 = 4'h4 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_492; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_685 = 4'h5 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_493; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_686 = 4'h6 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_494; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_687 = 4'h7 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_495; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_688 = 4'h8 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_496; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_689 = 4'h9 == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_497; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_690 = 4'ha == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_498; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_691 = 4'hb == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_499; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_692 = 4'hc == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_500; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_693 = 4'hd == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_501; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_694 = 4'he == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_502; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_695 = 4'hf == _full_T_4 ? _inst_queue_pc_T_5 : _GEN_503; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [1:0] _inst_queue_inst_T_6 = io_in_bits_offset + 2'h2; // @[IQueue.scala 55:74]
  wire [31:0] _GEN_713 = 2'h1 == _inst_queue_inst_T_6 ? in_inst_1 : in_inst_0; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_714 = 2'h2 == _inst_queue_inst_T_6 ? in_inst_2 : _GEN_713; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_715 = 2'h3 == _inst_queue_inst_T_6 ? in_inst_3 : _GEN_714; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_696 = 4'h0 == _full_T_4 ? _GEN_715 : _GEN_504; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_697 = 4'h1 == _full_T_4 ? _GEN_715 : _GEN_505; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_698 = 4'h2 == _full_T_4 ? _GEN_715 : _GEN_506; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_699 = 4'h3 == _full_T_4 ? _GEN_715 : _GEN_507; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_700 = 4'h4 == _full_T_4 ? _GEN_715 : _GEN_508; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_701 = 4'h5 == _full_T_4 ? _GEN_715 : _GEN_509; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_702 = 4'h6 == _full_T_4 ? _GEN_715 : _GEN_510; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_703 = 4'h7 == _full_T_4 ? _GEN_715 : _GEN_511; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_704 = 4'h8 == _full_T_4 ? _GEN_715 : _GEN_512; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_705 = 4'h9 == _full_T_4 ? _GEN_715 : _GEN_513; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_706 = 4'ha == _full_T_4 ? _GEN_715 : _GEN_514; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_707 = 4'hb == _full_T_4 ? _GEN_715 : _GEN_515; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_708 = 4'hc == _full_T_4 ? _GEN_715 : _GEN_516; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_709 = 4'hd == _full_T_4 ? _GEN_715 : _GEN_517; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_710 = 4'he == _full_T_4 ? _GEN_715 : _GEN_518; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_711 = 4'hf == _full_T_4 ? _GEN_715 : _GEN_519; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire  _GEN_716 = 4'h0 == _full_T_4 ? 1'h0 : _GEN_632; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_717 = 4'h1 == _full_T_4 ? 1'h0 : _GEN_633; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_718 = 4'h2 == _full_T_4 ? 1'h0 : _GEN_634; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_719 = 4'h3 == _full_T_4 ? 1'h0 : _GEN_635; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_720 = 4'h4 == _full_T_4 ? 1'h0 : _GEN_636; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_721 = 4'h5 == _full_T_4 ? 1'h0 : _GEN_637; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_722 = 4'h6 == _full_T_4 ? 1'h0 : _GEN_638; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_723 = 4'h7 == _full_T_4 ? 1'h0 : _GEN_639; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_724 = 4'h8 == _full_T_4 ? 1'h0 : _GEN_640; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_725 = 4'h9 == _full_T_4 ? 1'h0 : _GEN_641; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_726 = 4'ha == _full_T_4 ? 1'h0 : _GEN_642; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_727 = 4'hb == _full_T_4 ? 1'h0 : _GEN_643; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_728 = 4'hc == _full_T_4 ? 1'h0 : _GEN_644; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_729 = 4'hd == _full_T_4 ? 1'h0 : _GEN_645; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_730 = 4'he == _full_T_4 ? 1'h0 : _GEN_646; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_731 = 4'hf == _full_T_4 ? 1'h0 : _GEN_647; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire [31:0] _GEN_732 = 4'h0 == _full_T_4 ? 32'h0 : _GEN_648; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_733 = 4'h1 == _full_T_4 ? 32'h0 : _GEN_649; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_734 = 4'h2 == _full_T_4 ? 32'h0 : _GEN_650; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_735 = 4'h3 == _full_T_4 ? 32'h0 : _GEN_651; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_736 = 4'h4 == _full_T_4 ? 32'h0 : _GEN_652; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_737 = 4'h5 == _full_T_4 ? 32'h0 : _GEN_653; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_738 = 4'h6 == _full_T_4 ? 32'h0 : _GEN_654; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_739 = 4'h7 == _full_T_4 ? 32'h0 : _GEN_655; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_740 = 4'h8 == _full_T_4 ? 32'h0 : _GEN_656; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_741 = 4'h9 == _full_T_4 ? 32'h0 : _GEN_657; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_742 = 4'ha == _full_T_4 ? 32'h0 : _GEN_658; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_743 = 4'hb == _full_T_4 ? 32'h0 : _GEN_659; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_744 = 4'hc == _full_T_4 ? 32'h0 : _GEN_660; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_745 = 4'hd == _full_T_4 ? 32'h0 : _GEN_661; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_746 = 4'he == _full_T_4 ? 32'h0 : _GEN_662; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_747 = 4'hf == _full_T_4 ? 32'h0 : _GEN_663; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [1:0] _GEN_748 = 4'h0 == _full_T_4 ? 2'h0 : _GEN_664; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_749 = 4'h1 == _full_T_4 ? 2'h0 : _GEN_665; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_750 = 4'h2 == _full_T_4 ? 2'h0 : _GEN_666; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_751 = 4'h3 == _full_T_4 ? 2'h0 : _GEN_667; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_752 = 4'h4 == _full_T_4 ? 2'h0 : _GEN_668; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_753 = 4'h5 == _full_T_4 ? 2'h0 : _GEN_669; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_754 = 4'h6 == _full_T_4 ? 2'h0 : _GEN_670; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_755 = 4'h7 == _full_T_4 ? 2'h0 : _GEN_671; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_756 = 4'h8 == _full_T_4 ? 2'h0 : _GEN_672; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_757 = 4'h9 == _full_T_4 ? 2'h0 : _GEN_673; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_758 = 4'ha == _full_T_4 ? 2'h0 : _GEN_674; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_759 = 4'hb == _full_T_4 ? 2'h0 : _GEN_675; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_760 = 4'hc == _full_T_4 ? 2'h0 : _GEN_676; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_761 = 4'hd == _full_T_4 ? 2'h0 : _GEN_677; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_762 = 4'he == _full_T_4 ? 2'h0 : _GEN_678; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_763 = 4'hf == _full_T_4 ? 2'h0 : _GEN_679; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire  _GEN_764 = 4'h0 == _full_T_4 | _GEN_568; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_765 = 4'h1 == _full_T_4 | _GEN_569; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_766 = 4'h2 == _full_T_4 | _GEN_570; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_767 = 4'h3 == _full_T_4 | _GEN_571; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_768 = 4'h4 == _full_T_4 | _GEN_572; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_769 = 4'h5 == _full_T_4 | _GEN_573; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_770 = 4'h6 == _full_T_4 | _GEN_574; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_771 = 4'h7 == _full_T_4 | _GEN_575; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_772 = 4'h8 == _full_T_4 | _GEN_576; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_773 = 4'h9 == _full_T_4 | _GEN_577; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_774 = 4'ha == _full_T_4 | _GEN_578; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_775 = 4'hb == _full_T_4 | _GEN_579; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_776 = 4'hc == _full_T_4 | _GEN_580; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_777 = 4'hd == _full_T_4 | _GEN_581; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_778 = 4'he == _full_T_4 | _GEN_582; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_779 = 4'hf == _full_T_4 | _GEN_583; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire [31:0] _GEN_780 = 2'h2 <= count ? _GEN_680 : _GEN_488; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_781 = 2'h2 <= count ? _GEN_681 : _GEN_489; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_782 = 2'h2 <= count ? _GEN_682 : _GEN_490; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_783 = 2'h2 <= count ? _GEN_683 : _GEN_491; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_784 = 2'h2 <= count ? _GEN_684 : _GEN_492; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_785 = 2'h2 <= count ? _GEN_685 : _GEN_493; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_786 = 2'h2 <= count ? _GEN_686 : _GEN_494; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_787 = 2'h2 <= count ? _GEN_687 : _GEN_495; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_788 = 2'h2 <= count ? _GEN_688 : _GEN_496; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_789 = 2'h2 <= count ? _GEN_689 : _GEN_497; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_790 = 2'h2 <= count ? _GEN_690 : _GEN_498; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_791 = 2'h2 <= count ? _GEN_691 : _GEN_499; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_792 = 2'h2 <= count ? _GEN_692 : _GEN_500; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_793 = 2'h2 <= count ? _GEN_693 : _GEN_501; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_794 = 2'h2 <= count ? _GEN_694 : _GEN_502; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_795 = 2'h2 <= count ? _GEN_695 : _GEN_503; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_796 = 2'h2 <= count ? _GEN_696 : _GEN_504; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_797 = 2'h2 <= count ? _GEN_697 : _GEN_505; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_798 = 2'h2 <= count ? _GEN_698 : _GEN_506; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_799 = 2'h2 <= count ? _GEN_699 : _GEN_507; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_800 = 2'h2 <= count ? _GEN_700 : _GEN_508; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_801 = 2'h2 <= count ? _GEN_701 : _GEN_509; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_802 = 2'h2 <= count ? _GEN_702 : _GEN_510; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_803 = 2'h2 <= count ? _GEN_703 : _GEN_511; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_804 = 2'h2 <= count ? _GEN_704 : _GEN_512; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_805 = 2'h2 <= count ? _GEN_705 : _GEN_513; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_806 = 2'h2 <= count ? _GEN_706 : _GEN_514; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_807 = 2'h2 <= count ? _GEN_707 : _GEN_515; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_808 = 2'h2 <= count ? _GEN_708 : _GEN_516; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_809 = 2'h2 <= count ? _GEN_709 : _GEN_517; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_810 = 2'h2 <= count ? _GEN_710 : _GEN_518; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_811 = 2'h2 <= count ? _GEN_711 : _GEN_519; // @[IQueue.scala 53:29]
  wire  _GEN_812 = 2'h2 <= count ? _GEN_716 : _GEN_632; // @[IQueue.scala 53:29]
  wire  _GEN_813 = 2'h2 <= count ? _GEN_717 : _GEN_633; // @[IQueue.scala 53:29]
  wire  _GEN_814 = 2'h2 <= count ? _GEN_718 : _GEN_634; // @[IQueue.scala 53:29]
  wire  _GEN_815 = 2'h2 <= count ? _GEN_719 : _GEN_635; // @[IQueue.scala 53:29]
  wire  _GEN_816 = 2'h2 <= count ? _GEN_720 : _GEN_636; // @[IQueue.scala 53:29]
  wire  _GEN_817 = 2'h2 <= count ? _GEN_721 : _GEN_637; // @[IQueue.scala 53:29]
  wire  _GEN_818 = 2'h2 <= count ? _GEN_722 : _GEN_638; // @[IQueue.scala 53:29]
  wire  _GEN_819 = 2'h2 <= count ? _GEN_723 : _GEN_639; // @[IQueue.scala 53:29]
  wire  _GEN_820 = 2'h2 <= count ? _GEN_724 : _GEN_640; // @[IQueue.scala 53:29]
  wire  _GEN_821 = 2'h2 <= count ? _GEN_725 : _GEN_641; // @[IQueue.scala 53:29]
  wire  _GEN_822 = 2'h2 <= count ? _GEN_726 : _GEN_642; // @[IQueue.scala 53:29]
  wire  _GEN_823 = 2'h2 <= count ? _GEN_727 : _GEN_643; // @[IQueue.scala 53:29]
  wire  _GEN_824 = 2'h2 <= count ? _GEN_728 : _GEN_644; // @[IQueue.scala 53:29]
  wire  _GEN_825 = 2'h2 <= count ? _GEN_729 : _GEN_645; // @[IQueue.scala 53:29]
  wire  _GEN_826 = 2'h2 <= count ? _GEN_730 : _GEN_646; // @[IQueue.scala 53:29]
  wire  _GEN_827 = 2'h2 <= count ? _GEN_731 : _GEN_647; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_828 = 2'h2 <= count ? _GEN_732 : _GEN_648; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_829 = 2'h2 <= count ? _GEN_733 : _GEN_649; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_830 = 2'h2 <= count ? _GEN_734 : _GEN_650; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_831 = 2'h2 <= count ? _GEN_735 : _GEN_651; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_832 = 2'h2 <= count ? _GEN_736 : _GEN_652; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_833 = 2'h2 <= count ? _GEN_737 : _GEN_653; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_834 = 2'h2 <= count ? _GEN_738 : _GEN_654; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_835 = 2'h2 <= count ? _GEN_739 : _GEN_655; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_836 = 2'h2 <= count ? _GEN_740 : _GEN_656; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_837 = 2'h2 <= count ? _GEN_741 : _GEN_657; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_838 = 2'h2 <= count ? _GEN_742 : _GEN_658; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_839 = 2'h2 <= count ? _GEN_743 : _GEN_659; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_840 = 2'h2 <= count ? _GEN_744 : _GEN_660; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_841 = 2'h2 <= count ? _GEN_745 : _GEN_661; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_842 = 2'h2 <= count ? _GEN_746 : _GEN_662; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_843 = 2'h2 <= count ? _GEN_747 : _GEN_663; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_844 = 2'h2 <= count ? _GEN_748 : _GEN_664; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_845 = 2'h2 <= count ? _GEN_749 : _GEN_665; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_846 = 2'h2 <= count ? _GEN_750 : _GEN_666; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_847 = 2'h2 <= count ? _GEN_751 : _GEN_667; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_848 = 2'h2 <= count ? _GEN_752 : _GEN_668; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_849 = 2'h2 <= count ? _GEN_753 : _GEN_669; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_850 = 2'h2 <= count ? _GEN_754 : _GEN_670; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_851 = 2'h2 <= count ? _GEN_755 : _GEN_671; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_852 = 2'h2 <= count ? _GEN_756 : _GEN_672; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_853 = 2'h2 <= count ? _GEN_757 : _GEN_673; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_854 = 2'h2 <= count ? _GEN_758 : _GEN_674; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_855 = 2'h2 <= count ? _GEN_759 : _GEN_675; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_856 = 2'h2 <= count ? _GEN_760 : _GEN_676; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_857 = 2'h2 <= count ? _GEN_761 : _GEN_677; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_858 = 2'h2 <= count ? _GEN_762 : _GEN_678; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_859 = 2'h2 <= count ? _GEN_763 : _GEN_679; // @[IQueue.scala 53:29]
  wire  _GEN_860 = 2'h2 <= count ? _GEN_764 : _GEN_568; // @[IQueue.scala 53:29]
  wire  _GEN_861 = 2'h2 <= count ? _GEN_765 : _GEN_569; // @[IQueue.scala 53:29]
  wire  _GEN_862 = 2'h2 <= count ? _GEN_766 : _GEN_570; // @[IQueue.scala 53:29]
  wire  _GEN_863 = 2'h2 <= count ? _GEN_767 : _GEN_571; // @[IQueue.scala 53:29]
  wire  _GEN_864 = 2'h2 <= count ? _GEN_768 : _GEN_572; // @[IQueue.scala 53:29]
  wire  _GEN_865 = 2'h2 <= count ? _GEN_769 : _GEN_573; // @[IQueue.scala 53:29]
  wire  _GEN_866 = 2'h2 <= count ? _GEN_770 : _GEN_574; // @[IQueue.scala 53:29]
  wire  _GEN_867 = 2'h2 <= count ? _GEN_771 : _GEN_575; // @[IQueue.scala 53:29]
  wire  _GEN_868 = 2'h2 <= count ? _GEN_772 : _GEN_576; // @[IQueue.scala 53:29]
  wire  _GEN_869 = 2'h2 <= count ? _GEN_773 : _GEN_577; // @[IQueue.scala 53:29]
  wire  _GEN_870 = 2'h2 <= count ? _GEN_774 : _GEN_578; // @[IQueue.scala 53:29]
  wire  _GEN_871 = 2'h2 <= count ? _GEN_775 : _GEN_579; // @[IQueue.scala 53:29]
  wire  _GEN_872 = 2'h2 <= count ? _GEN_776 : _GEN_580; // @[IQueue.scala 53:29]
  wire  _GEN_873 = 2'h2 <= count ? _GEN_777 : _GEN_581; // @[IQueue.scala 53:29]
  wire  _GEN_874 = 2'h2 <= count ? _GEN_778 : _GEN_582; // @[IQueue.scala 53:29]
  wire  _GEN_875 = 2'h2 <= count ? _GEN_779 : _GEN_583; // @[IQueue.scala 53:29]
  wire  _GEN_876 = 4'h0 == _T_15 ? io_in_bits_bp_br_taken : _GEN_812; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_877 = 4'h1 == _T_15 ? io_in_bits_bp_br_taken : _GEN_813; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_878 = 4'h2 == _T_15 ? io_in_bits_bp_br_taken : _GEN_814; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_879 = 4'h3 == _T_15 ? io_in_bits_bp_br_taken : _GEN_815; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_880 = 4'h4 == _T_15 ? io_in_bits_bp_br_taken : _GEN_816; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_881 = 4'h5 == _T_15 ? io_in_bits_bp_br_taken : _GEN_817; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_882 = 4'h6 == _T_15 ? io_in_bits_bp_br_taken : _GEN_818; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_883 = 4'h7 == _T_15 ? io_in_bits_bp_br_taken : _GEN_819; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_884 = 4'h8 == _T_15 ? io_in_bits_bp_br_taken : _GEN_820; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_885 = 4'h9 == _T_15 ? io_in_bits_bp_br_taken : _GEN_821; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_886 = 4'ha == _T_15 ? io_in_bits_bp_br_taken : _GEN_822; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_887 = 4'hb == _T_15 ? io_in_bits_bp_br_taken : _GEN_823; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_888 = 4'hc == _T_15 ? io_in_bits_bp_br_taken : _GEN_824; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_889 = 4'hd == _T_15 ? io_in_bits_bp_br_taken : _GEN_825; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_890 = 4'he == _T_15 ? io_in_bits_bp_br_taken : _GEN_826; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_891 = 4'hf == _T_15 ? io_in_bits_bp_br_taken : _GEN_827; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire [31:0] _GEN_892 = 4'h0 == _T_15 ? io_in_bits_bp_br_target : _GEN_828; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_893 = 4'h1 == _T_15 ? io_in_bits_bp_br_target : _GEN_829; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_894 = 4'h2 == _T_15 ? io_in_bits_bp_br_target : _GEN_830; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_895 = 4'h3 == _T_15 ? io_in_bits_bp_br_target : _GEN_831; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_896 = 4'h4 == _T_15 ? io_in_bits_bp_br_target : _GEN_832; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_897 = 4'h5 == _T_15 ? io_in_bits_bp_br_target : _GEN_833; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_898 = 4'h6 == _T_15 ? io_in_bits_bp_br_target : _GEN_834; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_899 = 4'h7 == _T_15 ? io_in_bits_bp_br_target : _GEN_835; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_900 = 4'h8 == _T_15 ? io_in_bits_bp_br_target : _GEN_836; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_901 = 4'h9 == _T_15 ? io_in_bits_bp_br_target : _GEN_837; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_902 = 4'ha == _T_15 ? io_in_bits_bp_br_target : _GEN_838; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_903 = 4'hb == _T_15 ? io_in_bits_bp_br_target : _GEN_839; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_904 = 4'hc == _T_15 ? io_in_bits_bp_br_target : _GEN_840; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_905 = 4'hd == _T_15 ? io_in_bits_bp_br_target : _GEN_841; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_906 = 4'he == _T_15 ? io_in_bits_bp_br_target : _GEN_842; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_907 = 4'hf == _T_15 ? io_in_bits_bp_br_target : _GEN_843; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [1:0] _GEN_908 = 4'h0 == _T_15 ? io_in_bits_bp_br_type : _GEN_844; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_909 = 4'h1 == _T_15 ? io_in_bits_bp_br_type : _GEN_845; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_910 = 4'h2 == _T_15 ? io_in_bits_bp_br_type : _GEN_846; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_911 = 4'h3 == _T_15 ? io_in_bits_bp_br_type : _GEN_847; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_912 = 4'h4 == _T_15 ? io_in_bits_bp_br_type : _GEN_848; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_913 = 4'h5 == _T_15 ? io_in_bits_bp_br_type : _GEN_849; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_914 = 4'h6 == _T_15 ? io_in_bits_bp_br_type : _GEN_850; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_915 = 4'h7 == _T_15 ? io_in_bits_bp_br_type : _GEN_851; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_916 = 4'h8 == _T_15 ? io_in_bits_bp_br_type : _GEN_852; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_917 = 4'h9 == _T_15 ? io_in_bits_bp_br_type : _GEN_853; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_918 = 4'ha == _T_15 ? io_in_bits_bp_br_type : _GEN_854; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_919 = 4'hb == _T_15 ? io_in_bits_bp_br_type : _GEN_855; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_920 = 4'hc == _T_15 ? io_in_bits_bp_br_type : _GEN_856; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_921 = 4'hd == _T_15 ? io_in_bits_bp_br_type : _GEN_857; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_922 = 4'he == _T_15 ? io_in_bits_bp_br_type : _GEN_858; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_923 = 4'hf == _T_15 ? io_in_bits_bp_br_type : _GEN_859; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire  _GEN_924 = has_bp_taken ? _GEN_876 : _GEN_812; // @[IQueue.scala 61:29]
  wire  _GEN_925 = has_bp_taken ? _GEN_877 : _GEN_813; // @[IQueue.scala 61:29]
  wire  _GEN_926 = has_bp_taken ? _GEN_878 : _GEN_814; // @[IQueue.scala 61:29]
  wire  _GEN_927 = has_bp_taken ? _GEN_879 : _GEN_815; // @[IQueue.scala 61:29]
  wire  _GEN_928 = has_bp_taken ? _GEN_880 : _GEN_816; // @[IQueue.scala 61:29]
  wire  _GEN_929 = has_bp_taken ? _GEN_881 : _GEN_817; // @[IQueue.scala 61:29]
  wire  _GEN_930 = has_bp_taken ? _GEN_882 : _GEN_818; // @[IQueue.scala 61:29]
  wire  _GEN_931 = has_bp_taken ? _GEN_883 : _GEN_819; // @[IQueue.scala 61:29]
  wire  _GEN_932 = has_bp_taken ? _GEN_884 : _GEN_820; // @[IQueue.scala 61:29]
  wire  _GEN_933 = has_bp_taken ? _GEN_885 : _GEN_821; // @[IQueue.scala 61:29]
  wire  _GEN_934 = has_bp_taken ? _GEN_886 : _GEN_822; // @[IQueue.scala 61:29]
  wire  _GEN_935 = has_bp_taken ? _GEN_887 : _GEN_823; // @[IQueue.scala 61:29]
  wire  _GEN_936 = has_bp_taken ? _GEN_888 : _GEN_824; // @[IQueue.scala 61:29]
  wire  _GEN_937 = has_bp_taken ? _GEN_889 : _GEN_825; // @[IQueue.scala 61:29]
  wire  _GEN_938 = has_bp_taken ? _GEN_890 : _GEN_826; // @[IQueue.scala 61:29]
  wire  _GEN_939 = has_bp_taken ? _GEN_891 : _GEN_827; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_940 = has_bp_taken ? _GEN_892 : _GEN_828; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_941 = has_bp_taken ? _GEN_893 : _GEN_829; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_942 = has_bp_taken ? _GEN_894 : _GEN_830; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_943 = has_bp_taken ? _GEN_895 : _GEN_831; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_944 = has_bp_taken ? _GEN_896 : _GEN_832; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_945 = has_bp_taken ? _GEN_897 : _GEN_833; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_946 = has_bp_taken ? _GEN_898 : _GEN_834; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_947 = has_bp_taken ? _GEN_899 : _GEN_835; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_948 = has_bp_taken ? _GEN_900 : _GEN_836; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_949 = has_bp_taken ? _GEN_901 : _GEN_837; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_950 = has_bp_taken ? _GEN_902 : _GEN_838; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_951 = has_bp_taken ? _GEN_903 : _GEN_839; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_952 = has_bp_taken ? _GEN_904 : _GEN_840; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_953 = has_bp_taken ? _GEN_905 : _GEN_841; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_954 = has_bp_taken ? _GEN_906 : _GEN_842; // @[IQueue.scala 61:29]
  wire [31:0] _GEN_955 = has_bp_taken ? _GEN_907 : _GEN_843; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_956 = has_bp_taken ? _GEN_908 : _GEN_844; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_957 = has_bp_taken ? _GEN_909 : _GEN_845; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_958 = has_bp_taken ? _GEN_910 : _GEN_846; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_959 = has_bp_taken ? _GEN_911 : _GEN_847; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_960 = has_bp_taken ? _GEN_912 : _GEN_848; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_961 = has_bp_taken ? _GEN_913 : _GEN_849; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_962 = has_bp_taken ? _GEN_914 : _GEN_850; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_963 = has_bp_taken ? _GEN_915 : _GEN_851; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_964 = has_bp_taken ? _GEN_916 : _GEN_852; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_965 = has_bp_taken ? _GEN_917 : _GEN_853; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_966 = has_bp_taken ? _GEN_918 : _GEN_854; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_967 = has_bp_taken ? _GEN_919 : _GEN_855; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_968 = has_bp_taken ? _GEN_920 : _GEN_856; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_969 = has_bp_taken ? _GEN_921 : _GEN_857; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_970 = has_bp_taken ? _GEN_922 : _GEN_858; // @[IQueue.scala 61:29]
  wire [1:0] _GEN_971 = has_bp_taken ? _GEN_923 : _GEN_859; // @[IQueue.scala 61:29]
  wire [31:0] _inst_queue_pc_T_7 = io_in_bits_pc + 32'hc; // @[IQueue.scala 54:60]
  wire [31:0] _GEN_972 = 4'h0 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_780; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_973 = 4'h1 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_781; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_974 = 4'h2 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_782; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_975 = 4'h3 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_783; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_976 = 4'h4 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_784; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_977 = 4'h5 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_785; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_978 = 4'h6 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_786; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_979 = 4'h7 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_787; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_980 = 4'h8 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_788; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_981 = 4'h9 == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_789; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_982 = 4'ha == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_790; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_983 = 4'hb == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_791; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_984 = 4'hc == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_792; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_985 = 4'hd == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_793; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_986 = 4'he == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_794; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [31:0] _GEN_987 = 4'hf == _full_T_8 ? _inst_queue_pc_T_7 : _GEN_795; // @[IQueue.scala 54:43 IQueue.scala 54:43]
  wire [1:0] _inst_queue_inst_T_8 = io_in_bits_offset + 2'h3; // @[IQueue.scala 55:74]
  wire [31:0] _GEN_1005 = 2'h1 == _inst_queue_inst_T_8 ? in_inst_1 : in_inst_0; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_1006 = 2'h2 == _inst_queue_inst_T_8 ? in_inst_2 : _GEN_1005; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_1007 = 2'h3 == _inst_queue_inst_T_8 ? in_inst_3 : _GEN_1006; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_988 = 4'h0 == _full_T_8 ? _GEN_1007 : _GEN_796; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_989 = 4'h1 == _full_T_8 ? _GEN_1007 : _GEN_797; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_990 = 4'h2 == _full_T_8 ? _GEN_1007 : _GEN_798; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_991 = 4'h3 == _full_T_8 ? _GEN_1007 : _GEN_799; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_992 = 4'h4 == _full_T_8 ? _GEN_1007 : _GEN_800; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_993 = 4'h5 == _full_T_8 ? _GEN_1007 : _GEN_801; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_994 = 4'h6 == _full_T_8 ? _GEN_1007 : _GEN_802; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_995 = 4'h7 == _full_T_8 ? _GEN_1007 : _GEN_803; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_996 = 4'h8 == _full_T_8 ? _GEN_1007 : _GEN_804; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_997 = 4'h9 == _full_T_8 ? _GEN_1007 : _GEN_805; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_998 = 4'ha == _full_T_8 ? _GEN_1007 : _GEN_806; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_999 = 4'hb == _full_T_8 ? _GEN_1007 : _GEN_807; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_1000 = 4'hc == _full_T_8 ? _GEN_1007 : _GEN_808; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_1001 = 4'hd == _full_T_8 ? _GEN_1007 : _GEN_809; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_1002 = 4'he == _full_T_8 ? _GEN_1007 : _GEN_810; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire [31:0] _GEN_1003 = 4'hf == _full_T_8 ? _GEN_1007 : _GEN_811; // @[IQueue.scala 55:45 IQueue.scala 55:45]
  wire  _GEN_1008 = 4'h0 == _full_T_8 ? 1'h0 : _GEN_924; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1009 = 4'h1 == _full_T_8 ? 1'h0 : _GEN_925; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1010 = 4'h2 == _full_T_8 ? 1'h0 : _GEN_926; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1011 = 4'h3 == _full_T_8 ? 1'h0 : _GEN_927; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1012 = 4'h4 == _full_T_8 ? 1'h0 : _GEN_928; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1013 = 4'h5 == _full_T_8 ? 1'h0 : _GEN_929; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1014 = 4'h6 == _full_T_8 ? 1'h0 : _GEN_930; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1015 = 4'h7 == _full_T_8 ? 1'h0 : _GEN_931; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1016 = 4'h8 == _full_T_8 ? 1'h0 : _GEN_932; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1017 = 4'h9 == _full_T_8 ? 1'h0 : _GEN_933; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1018 = 4'ha == _full_T_8 ? 1'h0 : _GEN_934; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1019 = 4'hb == _full_T_8 ? 1'h0 : _GEN_935; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1020 = 4'hc == _full_T_8 ? 1'h0 : _GEN_936; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1021 = 4'hd == _full_T_8 ? 1'h0 : _GEN_937; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1022 = 4'he == _full_T_8 ? 1'h0 : _GEN_938; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire  _GEN_1023 = 4'hf == _full_T_8 ? 1'h0 : _GEN_939; // @[IQueue.scala 56:52 IQueue.scala 56:52]
  wire [31:0] _GEN_1024 = 4'h0 == _full_T_8 ? 32'h0 : _GEN_940; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1025 = 4'h1 == _full_T_8 ? 32'h0 : _GEN_941; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1026 = 4'h2 == _full_T_8 ? 32'h0 : _GEN_942; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1027 = 4'h3 == _full_T_8 ? 32'h0 : _GEN_943; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1028 = 4'h4 == _full_T_8 ? 32'h0 : _GEN_944; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1029 = 4'h5 == _full_T_8 ? 32'h0 : _GEN_945; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1030 = 4'h6 == _full_T_8 ? 32'h0 : _GEN_946; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1031 = 4'h7 == _full_T_8 ? 32'h0 : _GEN_947; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1032 = 4'h8 == _full_T_8 ? 32'h0 : _GEN_948; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1033 = 4'h9 == _full_T_8 ? 32'h0 : _GEN_949; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1034 = 4'ha == _full_T_8 ? 32'h0 : _GEN_950; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1035 = 4'hb == _full_T_8 ? 32'h0 : _GEN_951; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1036 = 4'hc == _full_T_8 ? 32'h0 : _GEN_952; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1037 = 4'hd == _full_T_8 ? 32'h0 : _GEN_953; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1038 = 4'he == _full_T_8 ? 32'h0 : _GEN_954; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [31:0] _GEN_1039 = 4'hf == _full_T_8 ? 32'h0 : _GEN_955; // @[IQueue.scala 57:53 IQueue.scala 57:53]
  wire [1:0] _GEN_1040 = 4'h0 == _full_T_8 ? 2'h0 : _GEN_956; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1041 = 4'h1 == _full_T_8 ? 2'h0 : _GEN_957; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1042 = 4'h2 == _full_T_8 ? 2'h0 : _GEN_958; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1043 = 4'h3 == _full_T_8 ? 2'h0 : _GEN_959; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1044 = 4'h4 == _full_T_8 ? 2'h0 : _GEN_960; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1045 = 4'h5 == _full_T_8 ? 2'h0 : _GEN_961; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1046 = 4'h6 == _full_T_8 ? 2'h0 : _GEN_962; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1047 = 4'h7 == _full_T_8 ? 2'h0 : _GEN_963; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1048 = 4'h8 == _full_T_8 ? 2'h0 : _GEN_964; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1049 = 4'h9 == _full_T_8 ? 2'h0 : _GEN_965; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1050 = 4'ha == _full_T_8 ? 2'h0 : _GEN_966; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1051 = 4'hb == _full_T_8 ? 2'h0 : _GEN_967; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1052 = 4'hc == _full_T_8 ? 2'h0 : _GEN_968; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1053 = 4'hd == _full_T_8 ? 2'h0 : _GEN_969; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1054 = 4'he == _full_T_8 ? 2'h0 : _GEN_970; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire [1:0] _GEN_1055 = 4'hf == _full_T_8 ? 2'h0 : _GEN_971; // @[IQueue.scala 58:51 IQueue.scala 58:51]
  wire  _GEN_1056 = 4'h0 == _full_T_8 | _GEN_860; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1057 = 4'h1 == _full_T_8 | _GEN_861; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1058 = 4'h2 == _full_T_8 | _GEN_862; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1059 = 4'h3 == _full_T_8 | _GEN_863; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1060 = 4'h4 == _full_T_8 | _GEN_864; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1061 = 4'h5 == _full_T_8 | _GEN_865; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1062 = 4'h6 == _full_T_8 | _GEN_866; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1063 = 4'h7 == _full_T_8 | _GEN_867; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1064 = 4'h8 == _full_T_8 | _GEN_868; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1065 = 4'h9 == _full_T_8 | _GEN_869; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1066 = 4'ha == _full_T_8 | _GEN_870; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1067 = 4'hb == _full_T_8 | _GEN_871; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1068 = 4'hc == _full_T_8 | _GEN_872; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1069 = 4'hd == _full_T_8 | _GEN_873; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1070 = 4'he == _full_T_8 | _GEN_874; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1071 = 4'hf == _full_T_8 | _GEN_875; // @[IQueue.scala 59:35 IQueue.scala 59:35]
  wire  _GEN_1104 = 2'h3 <= count ? _GEN_1008 : _GEN_924; // @[IQueue.scala 53:29]
  wire  _GEN_1105 = 2'h3 <= count ? _GEN_1009 : _GEN_925; // @[IQueue.scala 53:29]
  wire  _GEN_1106 = 2'h3 <= count ? _GEN_1010 : _GEN_926; // @[IQueue.scala 53:29]
  wire  _GEN_1107 = 2'h3 <= count ? _GEN_1011 : _GEN_927; // @[IQueue.scala 53:29]
  wire  _GEN_1108 = 2'h3 <= count ? _GEN_1012 : _GEN_928; // @[IQueue.scala 53:29]
  wire  _GEN_1109 = 2'h3 <= count ? _GEN_1013 : _GEN_929; // @[IQueue.scala 53:29]
  wire  _GEN_1110 = 2'h3 <= count ? _GEN_1014 : _GEN_930; // @[IQueue.scala 53:29]
  wire  _GEN_1111 = 2'h3 <= count ? _GEN_1015 : _GEN_931; // @[IQueue.scala 53:29]
  wire  _GEN_1112 = 2'h3 <= count ? _GEN_1016 : _GEN_932; // @[IQueue.scala 53:29]
  wire  _GEN_1113 = 2'h3 <= count ? _GEN_1017 : _GEN_933; // @[IQueue.scala 53:29]
  wire  _GEN_1114 = 2'h3 <= count ? _GEN_1018 : _GEN_934; // @[IQueue.scala 53:29]
  wire  _GEN_1115 = 2'h3 <= count ? _GEN_1019 : _GEN_935; // @[IQueue.scala 53:29]
  wire  _GEN_1116 = 2'h3 <= count ? _GEN_1020 : _GEN_936; // @[IQueue.scala 53:29]
  wire  _GEN_1117 = 2'h3 <= count ? _GEN_1021 : _GEN_937; // @[IQueue.scala 53:29]
  wire  _GEN_1118 = 2'h3 <= count ? _GEN_1022 : _GEN_938; // @[IQueue.scala 53:29]
  wire  _GEN_1119 = 2'h3 <= count ? _GEN_1023 : _GEN_939; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1120 = 2'h3 <= count ? _GEN_1024 : _GEN_940; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1121 = 2'h3 <= count ? _GEN_1025 : _GEN_941; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1122 = 2'h3 <= count ? _GEN_1026 : _GEN_942; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1123 = 2'h3 <= count ? _GEN_1027 : _GEN_943; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1124 = 2'h3 <= count ? _GEN_1028 : _GEN_944; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1125 = 2'h3 <= count ? _GEN_1029 : _GEN_945; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1126 = 2'h3 <= count ? _GEN_1030 : _GEN_946; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1127 = 2'h3 <= count ? _GEN_1031 : _GEN_947; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1128 = 2'h3 <= count ? _GEN_1032 : _GEN_948; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1129 = 2'h3 <= count ? _GEN_1033 : _GEN_949; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1130 = 2'h3 <= count ? _GEN_1034 : _GEN_950; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1131 = 2'h3 <= count ? _GEN_1035 : _GEN_951; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1132 = 2'h3 <= count ? _GEN_1036 : _GEN_952; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1133 = 2'h3 <= count ? _GEN_1037 : _GEN_953; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1134 = 2'h3 <= count ? _GEN_1038 : _GEN_954; // @[IQueue.scala 53:29]
  wire [31:0] _GEN_1135 = 2'h3 <= count ? _GEN_1039 : _GEN_955; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1136 = 2'h3 <= count ? _GEN_1040 : _GEN_956; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1137 = 2'h3 <= count ? _GEN_1041 : _GEN_957; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1138 = 2'h3 <= count ? _GEN_1042 : _GEN_958; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1139 = 2'h3 <= count ? _GEN_1043 : _GEN_959; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1140 = 2'h3 <= count ? _GEN_1044 : _GEN_960; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1141 = 2'h3 <= count ? _GEN_1045 : _GEN_961; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1142 = 2'h3 <= count ? _GEN_1046 : _GEN_962; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1143 = 2'h3 <= count ? _GEN_1047 : _GEN_963; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1144 = 2'h3 <= count ? _GEN_1048 : _GEN_964; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1145 = 2'h3 <= count ? _GEN_1049 : _GEN_965; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1146 = 2'h3 <= count ? _GEN_1050 : _GEN_966; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1147 = 2'h3 <= count ? _GEN_1051 : _GEN_967; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1148 = 2'h3 <= count ? _GEN_1052 : _GEN_968; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1149 = 2'h3 <= count ? _GEN_1053 : _GEN_969; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1150 = 2'h3 <= count ? _GEN_1054 : _GEN_970; // @[IQueue.scala 53:29]
  wire [1:0] _GEN_1151 = 2'h3 <= count ? _GEN_1055 : _GEN_971; // @[IQueue.scala 53:29]
  wire  _GEN_1152 = 2'h3 <= count ? _GEN_1056 : _GEN_860; // @[IQueue.scala 53:29]
  wire  _GEN_1153 = 2'h3 <= count ? _GEN_1057 : _GEN_861; // @[IQueue.scala 53:29]
  wire  _GEN_1154 = 2'h3 <= count ? _GEN_1058 : _GEN_862; // @[IQueue.scala 53:29]
  wire  _GEN_1155 = 2'h3 <= count ? _GEN_1059 : _GEN_863; // @[IQueue.scala 53:29]
  wire  _GEN_1156 = 2'h3 <= count ? _GEN_1060 : _GEN_864; // @[IQueue.scala 53:29]
  wire  _GEN_1157 = 2'h3 <= count ? _GEN_1061 : _GEN_865; // @[IQueue.scala 53:29]
  wire  _GEN_1158 = 2'h3 <= count ? _GEN_1062 : _GEN_866; // @[IQueue.scala 53:29]
  wire  _GEN_1159 = 2'h3 <= count ? _GEN_1063 : _GEN_867; // @[IQueue.scala 53:29]
  wire  _GEN_1160 = 2'h3 <= count ? _GEN_1064 : _GEN_868; // @[IQueue.scala 53:29]
  wire  _GEN_1161 = 2'h3 <= count ? _GEN_1065 : _GEN_869; // @[IQueue.scala 53:29]
  wire  _GEN_1162 = 2'h3 <= count ? _GEN_1066 : _GEN_870; // @[IQueue.scala 53:29]
  wire  _GEN_1163 = 2'h3 <= count ? _GEN_1067 : _GEN_871; // @[IQueue.scala 53:29]
  wire  _GEN_1164 = 2'h3 <= count ? _GEN_1068 : _GEN_872; // @[IQueue.scala 53:29]
  wire  _GEN_1165 = 2'h3 <= count ? _GEN_1069 : _GEN_873; // @[IQueue.scala 53:29]
  wire  _GEN_1166 = 2'h3 <= count ? _GEN_1070 : _GEN_874; // @[IQueue.scala 53:29]
  wire  _GEN_1167 = 2'h3 <= count ? _GEN_1071 : _GEN_875; // @[IQueue.scala 53:29]
  wire  _GEN_1168 = 4'h0 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1104; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1169 = 4'h1 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1105; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1170 = 4'h2 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1106; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1171 = 4'h3 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1107; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1172 = 4'h4 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1108; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1173 = 4'h5 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1109; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1174 = 4'h6 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1110; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1175 = 4'h7 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1111; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1176 = 4'h8 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1112; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1177 = 4'h9 == _T_15 ? io_in_bits_bp_br_taken : _GEN_1113; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1178 = 4'ha == _T_15 ? io_in_bits_bp_br_taken : _GEN_1114; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1179 = 4'hb == _T_15 ? io_in_bits_bp_br_taken : _GEN_1115; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1180 = 4'hc == _T_15 ? io_in_bits_bp_br_taken : _GEN_1116; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1181 = 4'hd == _T_15 ? io_in_bits_bp_br_taken : _GEN_1117; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1182 = 4'he == _T_15 ? io_in_bits_bp_br_taken : _GEN_1118; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire  _GEN_1183 = 4'hf == _T_15 ? io_in_bits_bp_br_taken : _GEN_1119; // @[IQueue.scala 62:54 IQueue.scala 62:54]
  wire [31:0] _GEN_1184 = 4'h0 == _T_15 ? io_in_bits_bp_br_target : _GEN_1120; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1185 = 4'h1 == _T_15 ? io_in_bits_bp_br_target : _GEN_1121; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1186 = 4'h2 == _T_15 ? io_in_bits_bp_br_target : _GEN_1122; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1187 = 4'h3 == _T_15 ? io_in_bits_bp_br_target : _GEN_1123; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1188 = 4'h4 == _T_15 ? io_in_bits_bp_br_target : _GEN_1124; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1189 = 4'h5 == _T_15 ? io_in_bits_bp_br_target : _GEN_1125; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1190 = 4'h6 == _T_15 ? io_in_bits_bp_br_target : _GEN_1126; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1191 = 4'h7 == _T_15 ? io_in_bits_bp_br_target : _GEN_1127; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1192 = 4'h8 == _T_15 ? io_in_bits_bp_br_target : _GEN_1128; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1193 = 4'h9 == _T_15 ? io_in_bits_bp_br_target : _GEN_1129; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1194 = 4'ha == _T_15 ? io_in_bits_bp_br_target : _GEN_1130; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1195 = 4'hb == _T_15 ? io_in_bits_bp_br_target : _GEN_1131; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1196 = 4'hc == _T_15 ? io_in_bits_bp_br_target : _GEN_1132; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1197 = 4'hd == _T_15 ? io_in_bits_bp_br_target : _GEN_1133; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1198 = 4'he == _T_15 ? io_in_bits_bp_br_target : _GEN_1134; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [31:0] _GEN_1199 = 4'hf == _T_15 ? io_in_bits_bp_br_target : _GEN_1135; // @[IQueue.scala 63:55 IQueue.scala 63:55]
  wire [1:0] _GEN_1200 = 4'h0 == _T_15 ? io_in_bits_bp_br_type : _GEN_1136; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1201 = 4'h1 == _T_15 ? io_in_bits_bp_br_type : _GEN_1137; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1202 = 4'h2 == _T_15 ? io_in_bits_bp_br_type : _GEN_1138; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1203 = 4'h3 == _T_15 ? io_in_bits_bp_br_type : _GEN_1139; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1204 = 4'h4 == _T_15 ? io_in_bits_bp_br_type : _GEN_1140; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1205 = 4'h5 == _T_15 ? io_in_bits_bp_br_type : _GEN_1141; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1206 = 4'h6 == _T_15 ? io_in_bits_bp_br_type : _GEN_1142; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1207 = 4'h7 == _T_15 ? io_in_bits_bp_br_type : _GEN_1143; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1208 = 4'h8 == _T_15 ? io_in_bits_bp_br_type : _GEN_1144; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1209 = 4'h9 == _T_15 ? io_in_bits_bp_br_type : _GEN_1145; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1210 = 4'ha == _T_15 ? io_in_bits_bp_br_type : _GEN_1146; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1211 = 4'hb == _T_15 ? io_in_bits_bp_br_type : _GEN_1147; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1212 = 4'hc == _T_15 ? io_in_bits_bp_br_type : _GEN_1148; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1213 = 4'hd == _T_15 ? io_in_bits_bp_br_type : _GEN_1149; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1214 = 4'he == _T_15 ? io_in_bits_bp_br_type : _GEN_1150; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire [1:0] _GEN_1215 = 4'hf == _T_15 ? io_in_bits_bp_br_type : _GEN_1151; // @[IQueue.scala 64:53 IQueue.scala 64:53]
  wire  _GEN_1344 = io_in_bits_uncache ? _GEN_80 : _GEN_1152; // @[IQueue.scala 43:31]
  wire  _GEN_1345 = io_in_bits_uncache ? _GEN_81 : _GEN_1153; // @[IQueue.scala 43:31]
  wire  _GEN_1346 = io_in_bits_uncache ? _GEN_82 : _GEN_1154; // @[IQueue.scala 43:31]
  wire  _GEN_1347 = io_in_bits_uncache ? _GEN_83 : _GEN_1155; // @[IQueue.scala 43:31]
  wire  _GEN_1348 = io_in_bits_uncache ? _GEN_84 : _GEN_1156; // @[IQueue.scala 43:31]
  wire  _GEN_1349 = io_in_bits_uncache ? _GEN_85 : _GEN_1157; // @[IQueue.scala 43:31]
  wire  _GEN_1350 = io_in_bits_uncache ? _GEN_86 : _GEN_1158; // @[IQueue.scala 43:31]
  wire  _GEN_1351 = io_in_bits_uncache ? _GEN_87 : _GEN_1159; // @[IQueue.scala 43:31]
  wire  _GEN_1352 = io_in_bits_uncache ? _GEN_88 : _GEN_1160; // @[IQueue.scala 43:31]
  wire  _GEN_1353 = io_in_bits_uncache ? _GEN_89 : _GEN_1161; // @[IQueue.scala 43:31]
  wire  _GEN_1354 = io_in_bits_uncache ? _GEN_90 : _GEN_1162; // @[IQueue.scala 43:31]
  wire  _GEN_1355 = io_in_bits_uncache ? _GEN_91 : _GEN_1163; // @[IQueue.scala 43:31]
  wire  _GEN_1356 = io_in_bits_uncache ? _GEN_92 : _GEN_1164; // @[IQueue.scala 43:31]
  wire  _GEN_1357 = io_in_bits_uncache ? _GEN_93 : _GEN_1165; // @[IQueue.scala 43:31]
  wire  _GEN_1358 = io_in_bits_uncache ? _GEN_94 : _GEN_1166; // @[IQueue.scala 43:31]
  wire  _GEN_1359 = io_in_bits_uncache ? _GEN_95 : _GEN_1167; // @[IQueue.scala 43:31]
  wire  _GEN_1441 = _T ? _GEN_1344 : valid_0; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1442 = _T ? _GEN_1345 : valid_1; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1443 = _T ? _GEN_1346 : valid_2; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1444 = _T ? _GEN_1347 : valid_3; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1445 = _T ? _GEN_1348 : valid_4; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1446 = _T ? _GEN_1349 : valid_5; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1447 = _T ? _GEN_1350 : valid_6; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1448 = _T ? _GEN_1351 : valid_7; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1449 = _T ? _GEN_1352 : valid_8; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1450 = _T ? _GEN_1353 : valid_9; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1451 = _T ? _GEN_1354 : valid_10; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1452 = _T ? _GEN_1355 : valid_11; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1453 = _T ? _GEN_1356 : valid_12; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1454 = _T ? _GEN_1357 : valid_13; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1455 = _T ? _GEN_1358 : valid_14; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _GEN_1456 = _T ? _GEN_1359 : valid_15; // @[IQueue.scala 42:21 IQueue.scala 26:22]
  wire  _T_77 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _out_counter_T_1 = out_counter + 4'h2; // @[IQueue.scala 73:34]
  wire [4:0] _T_78 = {{1'd0}, out_counter}; // @[IQueue.scala 75:27]
  wire  _GEN_1458 = 4'h0 == _T_78[3:0] ? 1'h0 : _GEN_1441; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1459 = 4'h1 == _T_78[3:0] ? 1'h0 : _GEN_1442; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1460 = 4'h2 == _T_78[3:0] ? 1'h0 : _GEN_1443; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1461 = 4'h3 == _T_78[3:0] ? 1'h0 : _GEN_1444; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1462 = 4'h4 == _T_78[3:0] ? 1'h0 : _GEN_1445; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1463 = 4'h5 == _T_78[3:0] ? 1'h0 : _GEN_1446; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1464 = 4'h6 == _T_78[3:0] ? 1'h0 : _GEN_1447; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1465 = 4'h7 == _T_78[3:0] ? 1'h0 : _GEN_1448; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1466 = 4'h8 == _T_78[3:0] ? 1'h0 : _GEN_1449; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1467 = 4'h9 == _T_78[3:0] ? 1'h0 : _GEN_1450; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1468 = 4'ha == _T_78[3:0] ? 1'h0 : _GEN_1451; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1469 = 4'hb == _T_78[3:0] ? 1'h0 : _GEN_1452; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1470 = 4'hc == _T_78[3:0] ? 1'h0 : _GEN_1453; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1471 = 4'hd == _T_78[3:0] ? 1'h0 : _GEN_1454; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1472 = 4'he == _T_78[3:0] ? 1'h0 : _GEN_1455; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1473 = 4'hf == _T_78[3:0] ? 1'h0 : _GEN_1456; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire [3:0] _T_81 = out_counter + 4'h1; // @[IQueue.scala 75:27]
  wire  _GEN_1474 = 4'h0 == _T_81 ? 1'h0 : _GEN_1458; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1475 = 4'h1 == _T_81 ? 1'h0 : _GEN_1459; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1476 = 4'h2 == _T_81 ? 1'h0 : _GEN_1460; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1477 = 4'h3 == _T_81 ? 1'h0 : _GEN_1461; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1478 = 4'h4 == _T_81 ? 1'h0 : _GEN_1462; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1479 = 4'h5 == _T_81 ? 1'h0 : _GEN_1463; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1480 = 4'h6 == _T_81 ? 1'h0 : _GEN_1464; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1481 = 4'h7 == _T_81 ? 1'h0 : _GEN_1465; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1482 = 4'h8 == _T_81 ? 1'h0 : _GEN_1466; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1483 = 4'h9 == _T_81 ? 1'h0 : _GEN_1467; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1484 = 4'ha == _T_81 ? 1'h0 : _GEN_1468; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1485 = 4'hb == _T_81 ? 1'h0 : _GEN_1469; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1486 = 4'hc == _T_81 ? 1'h0 : _GEN_1470; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1487 = 4'hd == _T_81 ? 1'h0 : _GEN_1471; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1488 = 4'he == _T_81 ? 1'h0 : _GEN_1472; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1489 = 4'hf == _T_81 ? 1'h0 : _GEN_1473; // @[IQueue.scala 75:34 IQueue.scala 75:34]
  wire  _GEN_1490 = 4'h0 == out_counter ? 1'h0 : _GEN_1441; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1491 = 4'h1 == out_counter ? 1'h0 : _GEN_1442; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1492 = 4'h2 == out_counter ? 1'h0 : _GEN_1443; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1493 = 4'h3 == out_counter ? 1'h0 : _GEN_1444; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1494 = 4'h4 == out_counter ? 1'h0 : _GEN_1445; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1495 = 4'h5 == out_counter ? 1'h0 : _GEN_1446; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1496 = 4'h6 == out_counter ? 1'h0 : _GEN_1447; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1497 = 4'h7 == out_counter ? 1'h0 : _GEN_1448; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1498 = 4'h8 == out_counter ? 1'h0 : _GEN_1449; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1499 = 4'h9 == out_counter ? 1'h0 : _GEN_1450; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1500 = 4'ha == out_counter ? 1'h0 : _GEN_1451; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1501 = 4'hb == out_counter ? 1'h0 : _GEN_1452; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1502 = 4'hc == out_counter ? 1'h0 : _GEN_1453; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1503 = 4'hd == out_counter ? 1'h0 : _GEN_1454; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1504 = 4'he == out_counter ? 1'h0 : _GEN_1455; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1505 = 4'hf == out_counter ? 1'h0 : _GEN_1456; // @[IQueue.scala 79:26 IQueue.scala 79:26]
  wire  _GEN_1541 = 4'h1 == _T_78[3:0] ? valid_1 : valid_0; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1542 = 4'h2 == _T_78[3:0] ? valid_2 : _GEN_1541; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1543 = 4'h3 == _T_78[3:0] ? valid_3 : _GEN_1542; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1544 = 4'h4 == _T_78[3:0] ? valid_4 : _GEN_1543; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1545 = 4'h5 == _T_78[3:0] ? valid_5 : _GEN_1544; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1546 = 4'h6 == _T_78[3:0] ? valid_6 : _GEN_1545; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1547 = 4'h7 == _T_78[3:0] ? valid_7 : _GEN_1546; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1548 = 4'h8 == _T_78[3:0] ? valid_8 : _GEN_1547; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1549 = 4'h9 == _T_78[3:0] ? valid_9 : _GEN_1548; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1550 = 4'ha == _T_78[3:0] ? valid_10 : _GEN_1549; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1551 = 4'hb == _T_78[3:0] ? valid_11 : _GEN_1550; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1552 = 4'hc == _T_78[3:0] ? valid_12 : _GEN_1551; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1553 = 4'hd == _T_78[3:0] ? valid_13 : _GEN_1552; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1554 = 4'he == _T_78[3:0] ? valid_14 : _GEN_1553; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire [31:0] _GEN_1557 = 4'h1 == _T_78[3:0] ? inst_queue_1_pc : inst_queue_0_pc; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1558 = 4'h2 == _T_78[3:0] ? inst_queue_2_pc : _GEN_1557; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1559 = 4'h3 == _T_78[3:0] ? inst_queue_3_pc : _GEN_1558; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1560 = 4'h4 == _T_78[3:0] ? inst_queue_4_pc : _GEN_1559; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1561 = 4'h5 == _T_78[3:0] ? inst_queue_5_pc : _GEN_1560; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1562 = 4'h6 == _T_78[3:0] ? inst_queue_6_pc : _GEN_1561; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1563 = 4'h7 == _T_78[3:0] ? inst_queue_7_pc : _GEN_1562; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1564 = 4'h8 == _T_78[3:0] ? inst_queue_8_pc : _GEN_1563; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1565 = 4'h9 == _T_78[3:0] ? inst_queue_9_pc : _GEN_1564; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1566 = 4'ha == _T_78[3:0] ? inst_queue_10_pc : _GEN_1565; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1567 = 4'hb == _T_78[3:0] ? inst_queue_11_pc : _GEN_1566; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1568 = 4'hc == _T_78[3:0] ? inst_queue_12_pc : _GEN_1567; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1569 = 4'hd == _T_78[3:0] ? inst_queue_13_pc : _GEN_1568; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1570 = 4'he == _T_78[3:0] ? inst_queue_14_pc : _GEN_1569; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1573 = 4'h1 == _T_78[3:0] ? inst_queue_1_inst : inst_queue_0_inst; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1574 = 4'h2 == _T_78[3:0] ? inst_queue_2_inst : _GEN_1573; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1575 = 4'h3 == _T_78[3:0] ? inst_queue_3_inst : _GEN_1574; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1576 = 4'h4 == _T_78[3:0] ? inst_queue_4_inst : _GEN_1575; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1577 = 4'h5 == _T_78[3:0] ? inst_queue_5_inst : _GEN_1576; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1578 = 4'h6 == _T_78[3:0] ? inst_queue_6_inst : _GEN_1577; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1579 = 4'h7 == _T_78[3:0] ? inst_queue_7_inst : _GEN_1578; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1580 = 4'h8 == _T_78[3:0] ? inst_queue_8_inst : _GEN_1579; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1581 = 4'h9 == _T_78[3:0] ? inst_queue_9_inst : _GEN_1580; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1582 = 4'ha == _T_78[3:0] ? inst_queue_10_inst : _GEN_1581; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1583 = 4'hb == _T_78[3:0] ? inst_queue_11_inst : _GEN_1582; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1584 = 4'hc == _T_78[3:0] ? inst_queue_12_inst : _GEN_1583; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1585 = 4'hd == _T_78[3:0] ? inst_queue_13_inst : _GEN_1584; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1586 = 4'he == _T_78[3:0] ? inst_queue_14_inst : _GEN_1585; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire  _GEN_1589 = 4'h1 == _T_78[3:0] ? inst_queue_1_bp_br_taken : inst_queue_0_bp_br_taken; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1590 = 4'h2 == _T_78[3:0] ? inst_queue_2_bp_br_taken : _GEN_1589; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1591 = 4'h3 == _T_78[3:0] ? inst_queue_3_bp_br_taken : _GEN_1590; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1592 = 4'h4 == _T_78[3:0] ? inst_queue_4_bp_br_taken : _GEN_1591; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1593 = 4'h5 == _T_78[3:0] ? inst_queue_5_bp_br_taken : _GEN_1592; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1594 = 4'h6 == _T_78[3:0] ? inst_queue_6_bp_br_taken : _GEN_1593; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1595 = 4'h7 == _T_78[3:0] ? inst_queue_7_bp_br_taken : _GEN_1594; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1596 = 4'h8 == _T_78[3:0] ? inst_queue_8_bp_br_taken : _GEN_1595; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1597 = 4'h9 == _T_78[3:0] ? inst_queue_9_bp_br_taken : _GEN_1596; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1598 = 4'ha == _T_78[3:0] ? inst_queue_10_bp_br_taken : _GEN_1597; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1599 = 4'hb == _T_78[3:0] ? inst_queue_11_bp_br_taken : _GEN_1598; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1600 = 4'hc == _T_78[3:0] ? inst_queue_12_bp_br_taken : _GEN_1599; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1601 = 4'hd == _T_78[3:0] ? inst_queue_13_bp_br_taken : _GEN_1600; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1602 = 4'he == _T_78[3:0] ? inst_queue_14_bp_br_taken : _GEN_1601; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire [31:0] _GEN_1605 = 4'h1 == _T_78[3:0] ? inst_queue_1_bp_br_target : inst_queue_0_bp_br_target; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1606 = 4'h2 == _T_78[3:0] ? inst_queue_2_bp_br_target : _GEN_1605; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1607 = 4'h3 == _T_78[3:0] ? inst_queue_3_bp_br_target : _GEN_1606; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1608 = 4'h4 == _T_78[3:0] ? inst_queue_4_bp_br_target : _GEN_1607; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1609 = 4'h5 == _T_78[3:0] ? inst_queue_5_bp_br_target : _GEN_1608; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1610 = 4'h6 == _T_78[3:0] ? inst_queue_6_bp_br_target : _GEN_1609; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1611 = 4'h7 == _T_78[3:0] ? inst_queue_7_bp_br_target : _GEN_1610; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1612 = 4'h8 == _T_78[3:0] ? inst_queue_8_bp_br_target : _GEN_1611; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1613 = 4'h9 == _T_78[3:0] ? inst_queue_9_bp_br_target : _GEN_1612; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1614 = 4'ha == _T_78[3:0] ? inst_queue_10_bp_br_target : _GEN_1613; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1615 = 4'hb == _T_78[3:0] ? inst_queue_11_bp_br_target : _GEN_1614; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1616 = 4'hc == _T_78[3:0] ? inst_queue_12_bp_br_target : _GEN_1615; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1617 = 4'hd == _T_78[3:0] ? inst_queue_13_bp_br_target : _GEN_1616; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1618 = 4'he == _T_78[3:0] ? inst_queue_14_bp_br_target : _GEN_1617; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [1:0] _GEN_1621 = 4'h1 == _T_78[3:0] ? inst_queue_1_bp_br_type : inst_queue_0_bp_br_type; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1622 = 4'h2 == _T_78[3:0] ? inst_queue_2_bp_br_type : _GEN_1621; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1623 = 4'h3 == _T_78[3:0] ? inst_queue_3_bp_br_type : _GEN_1622; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1624 = 4'h4 == _T_78[3:0] ? inst_queue_4_bp_br_type : _GEN_1623; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1625 = 4'h5 == _T_78[3:0] ? inst_queue_5_bp_br_type : _GEN_1624; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1626 = 4'h6 == _T_78[3:0] ? inst_queue_6_bp_br_type : _GEN_1625; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1627 = 4'h7 == _T_78[3:0] ? inst_queue_7_bp_br_type : _GEN_1626; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1628 = 4'h8 == _T_78[3:0] ? inst_queue_8_bp_br_type : _GEN_1627; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1629 = 4'h9 == _T_78[3:0] ? inst_queue_9_bp_br_type : _GEN_1628; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1630 = 4'ha == _T_78[3:0] ? inst_queue_10_bp_br_type : _GEN_1629; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1631 = 4'hb == _T_78[3:0] ? inst_queue_11_bp_br_type : _GEN_1630; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1632 = 4'hc == _T_78[3:0] ? inst_queue_12_bp_br_type : _GEN_1631; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1633 = 4'hd == _T_78[3:0] ? inst_queue_13_bp_br_type : _GEN_1632; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1634 = 4'he == _T_78[3:0] ? inst_queue_14_bp_br_type : _GEN_1633; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire  _GEN_1637 = 4'h1 == _T_81 ? valid_1 : valid_0; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1638 = 4'h2 == _T_81 ? valid_2 : _GEN_1637; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1639 = 4'h3 == _T_81 ? valid_3 : _GEN_1638; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1640 = 4'h4 == _T_81 ? valid_4 : _GEN_1639; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1641 = 4'h5 == _T_81 ? valid_5 : _GEN_1640; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1642 = 4'h6 == _T_81 ? valid_6 : _GEN_1641; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1643 = 4'h7 == _T_81 ? valid_7 : _GEN_1642; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1644 = 4'h8 == _T_81 ? valid_8 : _GEN_1643; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1645 = 4'h9 == _T_81 ? valid_9 : _GEN_1644; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1646 = 4'ha == _T_81 ? valid_10 : _GEN_1645; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1647 = 4'hb == _T_81 ? valid_11 : _GEN_1646; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1648 = 4'hc == _T_81 ? valid_12 : _GEN_1647; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1649 = 4'hd == _T_81 ? valid_13 : _GEN_1648; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire  _GEN_1650 = 4'he == _T_81 ? valid_14 : _GEN_1649; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  wire [31:0] _GEN_1653 = 4'h1 == _T_81 ? inst_queue_1_pc : inst_queue_0_pc; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1654 = 4'h2 == _T_81 ? inst_queue_2_pc : _GEN_1653; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1655 = 4'h3 == _T_81 ? inst_queue_3_pc : _GEN_1654; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1656 = 4'h4 == _T_81 ? inst_queue_4_pc : _GEN_1655; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1657 = 4'h5 == _T_81 ? inst_queue_5_pc : _GEN_1656; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1658 = 4'h6 == _T_81 ? inst_queue_6_pc : _GEN_1657; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1659 = 4'h7 == _T_81 ? inst_queue_7_pc : _GEN_1658; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1660 = 4'h8 == _T_81 ? inst_queue_8_pc : _GEN_1659; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1661 = 4'h9 == _T_81 ? inst_queue_9_pc : _GEN_1660; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1662 = 4'ha == _T_81 ? inst_queue_10_pc : _GEN_1661; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1663 = 4'hb == _T_81 ? inst_queue_11_pc : _GEN_1662; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1664 = 4'hc == _T_81 ? inst_queue_12_pc : _GEN_1663; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1665 = 4'hd == _T_81 ? inst_queue_13_pc : _GEN_1664; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1666 = 4'he == _T_81 ? inst_queue_14_pc : _GEN_1665; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  wire [31:0] _GEN_1669 = 4'h1 == _T_81 ? inst_queue_1_inst : inst_queue_0_inst; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1670 = 4'h2 == _T_81 ? inst_queue_2_inst : _GEN_1669; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1671 = 4'h3 == _T_81 ? inst_queue_3_inst : _GEN_1670; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1672 = 4'h4 == _T_81 ? inst_queue_4_inst : _GEN_1671; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1673 = 4'h5 == _T_81 ? inst_queue_5_inst : _GEN_1672; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1674 = 4'h6 == _T_81 ? inst_queue_6_inst : _GEN_1673; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1675 = 4'h7 == _T_81 ? inst_queue_7_inst : _GEN_1674; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1676 = 4'h8 == _T_81 ? inst_queue_8_inst : _GEN_1675; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1677 = 4'h9 == _T_81 ? inst_queue_9_inst : _GEN_1676; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1678 = 4'ha == _T_81 ? inst_queue_10_inst : _GEN_1677; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1679 = 4'hb == _T_81 ? inst_queue_11_inst : _GEN_1678; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1680 = 4'hc == _T_81 ? inst_queue_12_inst : _GEN_1679; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1681 = 4'hd == _T_81 ? inst_queue_13_inst : _GEN_1680; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire [31:0] _GEN_1682 = 4'he == _T_81 ? inst_queue_14_inst : _GEN_1681; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  wire  _GEN_1685 = 4'h1 == _T_81 ? inst_queue_1_bp_br_taken : inst_queue_0_bp_br_taken; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1686 = 4'h2 == _T_81 ? inst_queue_2_bp_br_taken : _GEN_1685; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1687 = 4'h3 == _T_81 ? inst_queue_3_bp_br_taken : _GEN_1686; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1688 = 4'h4 == _T_81 ? inst_queue_4_bp_br_taken : _GEN_1687; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1689 = 4'h5 == _T_81 ? inst_queue_5_bp_br_taken : _GEN_1688; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1690 = 4'h6 == _T_81 ? inst_queue_6_bp_br_taken : _GEN_1689; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1691 = 4'h7 == _T_81 ? inst_queue_7_bp_br_taken : _GEN_1690; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1692 = 4'h8 == _T_81 ? inst_queue_8_bp_br_taken : _GEN_1691; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1693 = 4'h9 == _T_81 ? inst_queue_9_bp_br_taken : _GEN_1692; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1694 = 4'ha == _T_81 ? inst_queue_10_bp_br_taken : _GEN_1693; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1695 = 4'hb == _T_81 ? inst_queue_11_bp_br_taken : _GEN_1694; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1696 = 4'hc == _T_81 ? inst_queue_12_bp_br_taken : _GEN_1695; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1697 = 4'hd == _T_81 ? inst_queue_13_bp_br_taken : _GEN_1696; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire  _GEN_1698 = 4'he == _T_81 ? inst_queue_14_bp_br_taken : _GEN_1697; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  wire [31:0] _GEN_1701 = 4'h1 == _T_81 ? inst_queue_1_bp_br_target : inst_queue_0_bp_br_target; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1702 = 4'h2 == _T_81 ? inst_queue_2_bp_br_target : _GEN_1701; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1703 = 4'h3 == _T_81 ? inst_queue_3_bp_br_target : _GEN_1702; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1704 = 4'h4 == _T_81 ? inst_queue_4_bp_br_target : _GEN_1703; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1705 = 4'h5 == _T_81 ? inst_queue_5_bp_br_target : _GEN_1704; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1706 = 4'h6 == _T_81 ? inst_queue_6_bp_br_target : _GEN_1705; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1707 = 4'h7 == _T_81 ? inst_queue_7_bp_br_target : _GEN_1706; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1708 = 4'h8 == _T_81 ? inst_queue_8_bp_br_target : _GEN_1707; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1709 = 4'h9 == _T_81 ? inst_queue_9_bp_br_target : _GEN_1708; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1710 = 4'ha == _T_81 ? inst_queue_10_bp_br_target : _GEN_1709; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1711 = 4'hb == _T_81 ? inst_queue_11_bp_br_target : _GEN_1710; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1712 = 4'hc == _T_81 ? inst_queue_12_bp_br_target : _GEN_1711; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1713 = 4'hd == _T_81 ? inst_queue_13_bp_br_target : _GEN_1712; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [31:0] _GEN_1714 = 4'he == _T_81 ? inst_queue_14_bp_br_target : _GEN_1713; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  wire [1:0] _GEN_1717 = 4'h1 == _T_81 ? inst_queue_1_bp_br_type : inst_queue_0_bp_br_type; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1718 = 4'h2 == _T_81 ? inst_queue_2_bp_br_type : _GEN_1717; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1719 = 4'h3 == _T_81 ? inst_queue_3_bp_br_type : _GEN_1718; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1720 = 4'h4 == _T_81 ? inst_queue_4_bp_br_type : _GEN_1719; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1721 = 4'h5 == _T_81 ? inst_queue_5_bp_br_type : _GEN_1720; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1722 = 4'h6 == _T_81 ? inst_queue_6_bp_br_type : _GEN_1721; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1723 = 4'h7 == _T_81 ? inst_queue_7_bp_br_type : _GEN_1722; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1724 = 4'h8 == _T_81 ? inst_queue_8_bp_br_type : _GEN_1723; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1725 = 4'h9 == _T_81 ? inst_queue_9_bp_br_type : _GEN_1724; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1726 = 4'ha == _T_81 ? inst_queue_10_bp_br_type : _GEN_1725; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1727 = 4'hb == _T_81 ? inst_queue_11_bp_br_type : _GEN_1726; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1728 = 4'hc == _T_81 ? inst_queue_12_bp_br_type : _GEN_1727; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1729 = 4'hd == _T_81 ? inst_queue_13_bp_br_type : _GEN_1728; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  wire [1:0] _GEN_1730 = 4'he == _T_81 ? inst_queue_14_bp_br_type : _GEN_1729; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  assign io_in_ready = ~full; // @[IQueue.scala 93:18]
  assign io_out_valid = ~frontend_reflush & io_out_bits_0_valid; // @[IQueue.scala 92:31]
  assign io_out_bits_0_valid = 4'hf == _T_78[3:0] ? valid_15 : _GEN_1554; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  assign io_out_bits_0_pc = 4'hf == _T_78[3:0] ? inst_queue_15_pc : _GEN_1570; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  assign io_out_bits_0_inst = 4'hf == _T_78[3:0] ? inst_queue_15_inst : _GEN_1586; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  assign io_out_bits_0_bp_br_taken = 4'hf == _T_78[3:0] ? inst_queue_15_bp_br_taken : _GEN_1602; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  assign io_out_bits_0_bp_br_target = 4'hf == _T_78[3:0] ? inst_queue_15_bp_br_target : _GEN_1618; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  assign io_out_bits_0_bp_br_type = 4'hf == _T_78[3:0] ? inst_queue_15_bp_br_type : _GEN_1634; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  assign io_out_bits_1_valid = 4'hf == _T_81 ? valid_15 : _GEN_1650; // @[IQueue.scala 84:26 IQueue.scala 84:26]
  assign io_out_bits_1_pc = 4'hf == _T_81 ? inst_queue_15_pc : _GEN_1666; // @[IQueue.scala 85:23 IQueue.scala 85:23]
  assign io_out_bits_1_inst = 4'hf == _T_81 ? inst_queue_15_inst : _GEN_1682; // @[IQueue.scala 86:25 IQueue.scala 86:25]
  assign io_out_bits_1_bp_br_taken = 4'hf == _T_81 ? inst_queue_15_bp_br_taken : _GEN_1698; // @[IQueue.scala 87:32 IQueue.scala 87:32]
  assign io_out_bits_1_bp_br_target = 4'hf == _T_81 ? inst_queue_15_bp_br_target : _GEN_1714; // @[IQueue.scala 88:33 IQueue.scala 88:33]
  assign io_out_bits_1_bp_br_type = 4'hf == _T_81 ? inst_queue_15_bp_br_type : _GEN_1730; // @[IQueue.scala 89:31 IQueue.scala 89:31]
  always @(posedge clock) begin
    if (reset) begin // @[IQueue.scala 22:27]
      in_counter <= 4'h0; // @[IQueue.scala 22:27]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      in_counter <= 4'h0; // @[IQueue.scala 97:16]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        in_counter <= _full_T_1; // @[IQueue.scala 50:18]
      end else begin
        in_counter <= _in_counter_T_5; // @[IQueue.scala 66:20]
      end
    end
    if (reset) begin // @[IQueue.scala 23:28]
      out_counter <= 4'h0; // @[IQueue.scala 23:28]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      out_counter <= 4'h0; // @[IQueue.scala 98:17]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        out_counter <= _out_counter_T_1; // @[IQueue.scala 73:19]
      end else begin
        out_counter <= _T_81; // @[IQueue.scala 78:19]
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_0_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h0 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_0_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_0_pc <= _GEN_972;
      end else begin
        inst_queue_0_pc <= _GEN_780;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_0_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h0 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_0_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_0_inst <= _GEN_988;
      end else begin
        inst_queue_0_inst <= _GEN_796;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_0_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h0 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_0_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_0_bp_br_taken <= _GEN_1168;
      end else begin
        inst_queue_0_bp_br_taken <= _GEN_1104;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_0_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h0 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_0_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_0_bp_br_target <= _GEN_1184;
      end else begin
        inst_queue_0_bp_br_target <= _GEN_1120;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_0_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h0 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_0_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_0_bp_br_type <= _GEN_1200;
      end else begin
        inst_queue_0_bp_br_type <= _GEN_1136;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_1_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h1 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_1_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_1_pc <= _GEN_973;
      end else begin
        inst_queue_1_pc <= _GEN_781;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_1_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h1 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_1_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_1_inst <= _GEN_989;
      end else begin
        inst_queue_1_inst <= _GEN_797;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_1_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h1 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_1_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_1_bp_br_taken <= _GEN_1169;
      end else begin
        inst_queue_1_bp_br_taken <= _GEN_1105;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_1_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h1 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_1_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_1_bp_br_target <= _GEN_1185;
      end else begin
        inst_queue_1_bp_br_target <= _GEN_1121;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_1_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h1 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_1_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_1_bp_br_type <= _GEN_1201;
      end else begin
        inst_queue_1_bp_br_type <= _GEN_1137;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_2_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h2 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_2_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_2_pc <= _GEN_974;
      end else begin
        inst_queue_2_pc <= _GEN_782;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_2_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h2 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_2_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_2_inst <= _GEN_990;
      end else begin
        inst_queue_2_inst <= _GEN_798;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_2_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h2 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_2_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_2_bp_br_taken <= _GEN_1170;
      end else begin
        inst_queue_2_bp_br_taken <= _GEN_1106;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_2_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h2 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_2_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_2_bp_br_target <= _GEN_1186;
      end else begin
        inst_queue_2_bp_br_target <= _GEN_1122;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_2_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h2 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_2_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_2_bp_br_type <= _GEN_1202;
      end else begin
        inst_queue_2_bp_br_type <= _GEN_1138;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_3_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h3 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_3_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_3_pc <= _GEN_975;
      end else begin
        inst_queue_3_pc <= _GEN_783;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_3_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h3 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_3_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_3_inst <= _GEN_991;
      end else begin
        inst_queue_3_inst <= _GEN_799;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_3_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h3 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_3_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_3_bp_br_taken <= _GEN_1171;
      end else begin
        inst_queue_3_bp_br_taken <= _GEN_1107;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_3_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h3 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_3_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_3_bp_br_target <= _GEN_1187;
      end else begin
        inst_queue_3_bp_br_target <= _GEN_1123;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_3_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h3 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_3_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_3_bp_br_type <= _GEN_1203;
      end else begin
        inst_queue_3_bp_br_type <= _GEN_1139;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_4_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h4 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_4_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_4_pc <= _GEN_976;
      end else begin
        inst_queue_4_pc <= _GEN_784;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_4_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h4 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_4_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_4_inst <= _GEN_992;
      end else begin
        inst_queue_4_inst <= _GEN_800;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_4_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h4 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_4_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_4_bp_br_taken <= _GEN_1172;
      end else begin
        inst_queue_4_bp_br_taken <= _GEN_1108;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_4_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h4 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_4_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_4_bp_br_target <= _GEN_1188;
      end else begin
        inst_queue_4_bp_br_target <= _GEN_1124;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_4_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h4 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_4_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_4_bp_br_type <= _GEN_1204;
      end else begin
        inst_queue_4_bp_br_type <= _GEN_1140;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_5_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h5 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_5_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_5_pc <= _GEN_977;
      end else begin
        inst_queue_5_pc <= _GEN_785;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_5_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h5 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_5_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_5_inst <= _GEN_993;
      end else begin
        inst_queue_5_inst <= _GEN_801;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_5_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h5 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_5_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_5_bp_br_taken <= _GEN_1173;
      end else begin
        inst_queue_5_bp_br_taken <= _GEN_1109;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_5_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h5 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_5_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_5_bp_br_target <= _GEN_1189;
      end else begin
        inst_queue_5_bp_br_target <= _GEN_1125;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_5_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h5 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_5_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_5_bp_br_type <= _GEN_1205;
      end else begin
        inst_queue_5_bp_br_type <= _GEN_1141;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_6_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h6 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_6_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_6_pc <= _GEN_978;
      end else begin
        inst_queue_6_pc <= _GEN_786;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_6_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h6 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_6_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_6_inst <= _GEN_994;
      end else begin
        inst_queue_6_inst <= _GEN_802;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_6_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h6 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_6_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_6_bp_br_taken <= _GEN_1174;
      end else begin
        inst_queue_6_bp_br_taken <= _GEN_1110;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_6_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h6 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_6_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_6_bp_br_target <= _GEN_1190;
      end else begin
        inst_queue_6_bp_br_target <= _GEN_1126;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_6_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h6 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_6_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_6_bp_br_type <= _GEN_1206;
      end else begin
        inst_queue_6_bp_br_type <= _GEN_1142;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_7_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h7 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_7_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_7_pc <= _GEN_979;
      end else begin
        inst_queue_7_pc <= _GEN_787;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_7_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h7 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_7_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_7_inst <= _GEN_995;
      end else begin
        inst_queue_7_inst <= _GEN_803;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_7_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h7 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_7_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_7_bp_br_taken <= _GEN_1175;
      end else begin
        inst_queue_7_bp_br_taken <= _GEN_1111;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_7_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h7 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_7_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_7_bp_br_target <= _GEN_1191;
      end else begin
        inst_queue_7_bp_br_target <= _GEN_1127;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_7_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h7 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_7_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_7_bp_br_type <= _GEN_1207;
      end else begin
        inst_queue_7_bp_br_type <= _GEN_1143;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_8_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h8 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_8_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_8_pc <= _GEN_980;
      end else begin
        inst_queue_8_pc <= _GEN_788;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_8_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h8 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_8_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_8_inst <= _GEN_996;
      end else begin
        inst_queue_8_inst <= _GEN_804;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_8_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h8 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_8_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_8_bp_br_taken <= _GEN_1176;
      end else begin
        inst_queue_8_bp_br_taken <= _GEN_1112;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_8_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h8 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_8_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_8_bp_br_target <= _GEN_1192;
      end else begin
        inst_queue_8_bp_br_target <= _GEN_1128;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_8_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h8 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_8_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_8_bp_br_type <= _GEN_1208;
      end else begin
        inst_queue_8_bp_br_type <= _GEN_1144;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_9_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h9 == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_9_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_9_pc <= _GEN_981;
      end else begin
        inst_queue_9_pc <= _GEN_789;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_9_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h9 == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_9_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_9_inst <= _GEN_997;
      end else begin
        inst_queue_9_inst <= _GEN_805;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_9_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h9 == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_9_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_9_bp_br_taken <= _GEN_1177;
      end else begin
        inst_queue_9_bp_br_taken <= _GEN_1113;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_9_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h9 == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_9_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_9_bp_br_target <= _GEN_1193;
      end else begin
        inst_queue_9_bp_br_target <= _GEN_1129;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_9_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'h9 == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_9_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_9_bp_br_type <= _GEN_1209;
      end else begin
        inst_queue_9_bp_br_type <= _GEN_1145;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_10_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'ha == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_10_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_10_pc <= _GEN_982;
      end else begin
        inst_queue_10_pc <= _GEN_790;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_10_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'ha == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_10_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_10_inst <= _GEN_998;
      end else begin
        inst_queue_10_inst <= _GEN_806;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_10_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'ha == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_10_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_10_bp_br_taken <= _GEN_1178;
      end else begin
        inst_queue_10_bp_br_taken <= _GEN_1114;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_10_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'ha == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_10_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_10_bp_br_target <= _GEN_1194;
      end else begin
        inst_queue_10_bp_br_target <= _GEN_1130;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_10_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'ha == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_10_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_10_bp_br_type <= _GEN_1210;
      end else begin
        inst_queue_10_bp_br_type <= _GEN_1146;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_11_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hb == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_11_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_11_pc <= _GEN_983;
      end else begin
        inst_queue_11_pc <= _GEN_791;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_11_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hb == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_11_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_11_inst <= _GEN_999;
      end else begin
        inst_queue_11_inst <= _GEN_807;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_11_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hb == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_11_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_11_bp_br_taken <= _GEN_1179;
      end else begin
        inst_queue_11_bp_br_taken <= _GEN_1115;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_11_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hb == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_11_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_11_bp_br_target <= _GEN_1195;
      end else begin
        inst_queue_11_bp_br_target <= _GEN_1131;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_11_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hb == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_11_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_11_bp_br_type <= _GEN_1211;
      end else begin
        inst_queue_11_bp_br_type <= _GEN_1147;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_12_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hc == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_12_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_12_pc <= _GEN_984;
      end else begin
        inst_queue_12_pc <= _GEN_792;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_12_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hc == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_12_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_12_inst <= _GEN_1000;
      end else begin
        inst_queue_12_inst <= _GEN_808;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_12_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hc == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_12_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_12_bp_br_taken <= _GEN_1180;
      end else begin
        inst_queue_12_bp_br_taken <= _GEN_1116;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_12_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hc == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_12_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_12_bp_br_target <= _GEN_1196;
      end else begin
        inst_queue_12_bp_br_target <= _GEN_1132;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_12_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hc == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_12_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_12_bp_br_type <= _GEN_1212;
      end else begin
        inst_queue_12_bp_br_type <= _GEN_1148;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_13_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hd == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_13_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_13_pc <= _GEN_985;
      end else begin
        inst_queue_13_pc <= _GEN_793;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_13_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hd == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_13_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_13_inst <= _GEN_1001;
      end else begin
        inst_queue_13_inst <= _GEN_809;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_13_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hd == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_13_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_13_bp_br_taken <= _GEN_1181;
      end else begin
        inst_queue_13_bp_br_taken <= _GEN_1117;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_13_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hd == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_13_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_13_bp_br_target <= _GEN_1197;
      end else begin
        inst_queue_13_bp_br_target <= _GEN_1133;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_13_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hd == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_13_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_13_bp_br_type <= _GEN_1213;
      end else begin
        inst_queue_13_bp_br_type <= _GEN_1149;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_14_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'he == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_14_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_14_pc <= _GEN_986;
      end else begin
        inst_queue_14_pc <= _GEN_794;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_14_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'he == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_14_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_14_inst <= _GEN_1002;
      end else begin
        inst_queue_14_inst <= _GEN_810;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_14_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'he == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_14_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_14_bp_br_taken <= _GEN_1182;
      end else begin
        inst_queue_14_bp_br_taken <= _GEN_1118;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_14_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'he == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_14_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_14_bp_br_target <= _GEN_1198;
      end else begin
        inst_queue_14_bp_br_target <= _GEN_1134;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_14_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'he == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_14_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_14_bp_br_type <= _GEN_1214;
      end else begin
        inst_queue_14_bp_br_type <= _GEN_1150;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_15_pc <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hf == in_counter) begin // @[IQueue.scala 44:33]
          inst_queue_15_pc <= io_in_bits_pc; // @[IQueue.scala 44:33]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_15_pc <= _GEN_987;
      end else begin
        inst_queue_15_pc <= _GEN_795;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_15_inst <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hf == in_counter) begin // @[IQueue.scala 45:35]
          inst_queue_15_inst <= in_inst_0; // @[IQueue.scala 45:35]
        end
      end else if (2'h3 <= count) begin // @[IQueue.scala 53:29]
        inst_queue_15_inst <= _GEN_1003;
      end else begin
        inst_queue_15_inst <= _GEN_811;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_15_bp_br_taken <= 1'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hf == in_counter) begin // @[IQueue.scala 46:42]
          inst_queue_15_bp_br_taken <= io_in_bits_bp_br_taken; // @[IQueue.scala 46:42]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_15_bp_br_taken <= _GEN_1183;
      end else begin
        inst_queue_15_bp_br_taken <= _GEN_1119;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_15_bp_br_target <= 32'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hf == in_counter) begin // @[IQueue.scala 47:43]
          inst_queue_15_bp_br_target <= io_in_bits_bp_br_target; // @[IQueue.scala 47:43]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_15_bp_br_target <= _GEN_1199;
      end else begin
        inst_queue_15_bp_br_target <= _GEN_1135;
      end
    end
    if (reset) begin // @[IQueue.scala 24:27]
      inst_queue_15_bp_br_type <= 2'h0; // @[IQueue.scala 24:27]
    end else if (_T) begin // @[IQueue.scala 42:21]
      if (io_in_bits_uncache) begin // @[IQueue.scala 43:31]
        if (4'hf == in_counter) begin // @[IQueue.scala 48:41]
          inst_queue_15_bp_br_type <= io_in_bits_bp_br_type; // @[IQueue.scala 48:41]
        end
      end else if (has_bp_taken) begin // @[IQueue.scala 61:29]
        inst_queue_15_bp_br_type <= _GEN_1215;
      end else begin
        inst_queue_15_bp_br_type <= _GEN_1151;
      end
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_0 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_0 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_0 <= _GEN_1474;
      end else begin
        valid_0 <= _GEN_1490;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_0 <= _GEN_1344;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_1 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_1 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_1 <= _GEN_1475;
      end else begin
        valid_1 <= _GEN_1491;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_1 <= _GEN_1345;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_2 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_2 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_2 <= _GEN_1476;
      end else begin
        valid_2 <= _GEN_1492;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_2 <= _GEN_1346;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_3 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_3 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_3 <= _GEN_1477;
      end else begin
        valid_3 <= _GEN_1493;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_3 <= _GEN_1347;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_4 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_4 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_4 <= _GEN_1478;
      end else begin
        valid_4 <= _GEN_1494;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_4 <= _GEN_1348;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_5 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_5 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_5 <= _GEN_1479;
      end else begin
        valid_5 <= _GEN_1495;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_5 <= _GEN_1349;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_6 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_6 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_6 <= _GEN_1480;
      end else begin
        valid_6 <= _GEN_1496;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_6 <= _GEN_1350;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_7 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_7 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_7 <= _GEN_1481;
      end else begin
        valid_7 <= _GEN_1497;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_7 <= _GEN_1351;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_8 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_8 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_8 <= _GEN_1482;
      end else begin
        valid_8 <= _GEN_1498;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_8 <= _GEN_1352;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_9 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_9 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_9 <= _GEN_1483;
      end else begin
        valid_9 <= _GEN_1499;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_9 <= _GEN_1353;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_10 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_10 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_10 <= _GEN_1484;
      end else begin
        valid_10 <= _GEN_1500;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_10 <= _GEN_1354;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_11 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_11 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_11 <= _GEN_1485;
      end else begin
        valid_11 <= _GEN_1501;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_11 <= _GEN_1355;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_12 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_12 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_12 <= _GEN_1486;
      end else begin
        valid_12 <= _GEN_1502;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_12 <= _GEN_1356;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_13 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_13 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_13 <= _GEN_1487;
      end else begin
        valid_13 <= _GEN_1503;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_13 <= _GEN_1357;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_14 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_14 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_14 <= _GEN_1488;
      end else begin
        valid_14 <= _GEN_1504;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_14 <= _GEN_1358;
    end
    if (reset) begin // @[IQueue.scala 26:22]
      valid_15 <= 1'h0; // @[IQueue.scala 26:22]
    end else if (reset | frontend_reflush) begin // @[IQueue.scala 96:37]
      valid_15 <= 1'h0; // @[IQueue.scala 100:16]
    end else if (_T_77) begin // @[IQueue.scala 71:22]
      if (io_out_bits_1_valid) begin // @[IQueue.scala 72:33]
        valid_15 <= _GEN_1489;
      end else begin
        valid_15 <= _GEN_1505;
      end
    end else if (_T) begin // @[IQueue.scala 42:21]
      valid_15 <= _GEN_1359;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_counter = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  out_counter = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  inst_queue_0_pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  inst_queue_0_inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  inst_queue_0_bp_br_taken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  inst_queue_0_bp_br_target = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  inst_queue_0_bp_br_type = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  inst_queue_1_pc = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  inst_queue_1_inst = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inst_queue_1_bp_br_taken = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  inst_queue_1_bp_br_target = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  inst_queue_1_bp_br_type = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  inst_queue_2_pc = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  inst_queue_2_inst = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  inst_queue_2_bp_br_taken = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inst_queue_2_bp_br_target = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  inst_queue_2_bp_br_type = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  inst_queue_3_pc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  inst_queue_3_inst = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  inst_queue_3_bp_br_taken = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inst_queue_3_bp_br_target = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  inst_queue_3_bp_br_type = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  inst_queue_4_pc = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  inst_queue_4_inst = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  inst_queue_4_bp_br_taken = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  inst_queue_4_bp_br_target = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  inst_queue_4_bp_br_type = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  inst_queue_5_pc = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  inst_queue_5_inst = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  inst_queue_5_bp_br_taken = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  inst_queue_5_bp_br_target = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  inst_queue_5_bp_br_type = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  inst_queue_6_pc = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  inst_queue_6_inst = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  inst_queue_6_bp_br_taken = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  inst_queue_6_bp_br_target = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  inst_queue_6_bp_br_type = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  inst_queue_7_pc = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  inst_queue_7_inst = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  inst_queue_7_bp_br_taken = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  inst_queue_7_bp_br_target = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  inst_queue_7_bp_br_type = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  inst_queue_8_pc = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  inst_queue_8_inst = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  inst_queue_8_bp_br_taken = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  inst_queue_8_bp_br_target = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  inst_queue_8_bp_br_type = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  inst_queue_9_pc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  inst_queue_9_inst = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  inst_queue_9_bp_br_taken = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  inst_queue_9_bp_br_target = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  inst_queue_9_bp_br_type = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  inst_queue_10_pc = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  inst_queue_10_inst = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  inst_queue_10_bp_br_taken = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  inst_queue_10_bp_br_target = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  inst_queue_10_bp_br_type = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  inst_queue_11_pc = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  inst_queue_11_inst = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  inst_queue_11_bp_br_taken = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  inst_queue_11_bp_br_target = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  inst_queue_11_bp_br_type = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  inst_queue_12_pc = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  inst_queue_12_inst = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  inst_queue_12_bp_br_taken = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  inst_queue_12_bp_br_target = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  inst_queue_12_bp_br_type = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  inst_queue_13_pc = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  inst_queue_13_inst = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  inst_queue_13_bp_br_taken = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  inst_queue_13_bp_br_target = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  inst_queue_13_bp_br_type = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  inst_queue_14_pc = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  inst_queue_14_inst = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  inst_queue_14_bp_br_taken = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  inst_queue_14_bp_br_target = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  inst_queue_14_bp_br_type = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  inst_queue_15_pc = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  inst_queue_15_inst = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  inst_queue_15_bp_br_taken = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  inst_queue_15_bp_br_target = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  inst_queue_15_bp_br_type = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  valid_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_1 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_2 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_3 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_4 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_5 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_6 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_7 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_8 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_9 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_10 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_11 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_12 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_13 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_14 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_15 = _RAND_97[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode_Entry(
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input         io_in_bp_br_taken,
  input  [31:0] io_in_bp_br_target,
  input  [1:0]  io_in_bp_br_type,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output [1:0]  io_out_src1,
  output [1:0]  io_out_src2,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_dest,
  output [63:0] io_out_imm,
  output [2:0]  io_out_fu_type,
  output [3:0]  io_out_bru_op,
  output [4:0]  io_out_alu_op,
  output [3:0]  io_out_lsu_op,
  output [2:0]  io_out_csr_op,
  output [3:0]  io_out_mdu_op,
  output        io_out_wen,
  output        io_out_rv64,
  output        io_out_bp_br_taken,
  output [31:0] io_out_bp_br_target,
  output [1:0]  io_out_bp_br_type
);
  wire [51:0] imm_i_hi = io_in_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [11:0] imm_i_lo = io_in_inst[31:20]; // @[IDU.scala 20:43]
  wire [63:0] imm_i = {imm_i_hi,imm_i_lo}; // @[Cat.scala 30:58]
  wire [6:0] imm_s_hi_lo = io_in_inst[31:25]; // @[IDU.scala 21:43]
  wire [4:0] imm_s_lo = io_in_inst[11:7]; // @[IDU.scala 21:57]
  wire [63:0] imm_s = {imm_i_hi,imm_s_hi_lo,imm_s_lo}; // @[Cat.scala 30:58]
  wire  imm_b_hi_hi_lo = io_in_inst[7]; // @[IDU.scala 22:43]
  wire [5:0] imm_b_hi_lo = io_in_inst[30:25]; // @[IDU.scala 22:52]
  wire [3:0] imm_b_lo_hi = io_in_inst[11:8]; // @[IDU.scala 22:66]
  wire [63:0] imm_b = {imm_i_hi,imm_b_hi_hi_lo,imm_b_hi_lo,imm_b_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_u_hi_hi = io_in_inst[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [19:0] imm_u_hi_lo = io_in_inst[31:12]; // @[IDU.scala 23:43]
  wire [63:0] imm_u = {imm_u_hi_hi,imm_u_hi_lo,12'h0}; // @[Cat.scala 30:58]
  wire [43:0] imm_j_hi_hi_hi = io_in_inst[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 72:12]
  wire [7:0] imm_j_hi_hi_lo = io_in_inst[19:12]; // @[IDU.scala 24:43]
  wire  imm_j_hi_lo = io_in_inst[20]; // @[IDU.scala 24:57]
  wire [9:0] imm_j_lo_hi = io_in_inst[30:21]; // @[IDU.scala 24:67]
  wire [63:0] imm_j = {imm_j_hi_hi_hi,imm_j_hi_hi_lo,imm_j_hi_lo,imm_j_lo_hi,1'h0}; // @[Cat.scala 30:58]
  wire [31:0] _information_T = io_in_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _information_T_1 = 32'h37 == _information_T; // @[Lookup.scala 31:38]
  wire  _information_T_3 = 32'h17 == _information_T; // @[Lookup.scala 31:38]
  wire  _information_T_5 = 32'h6f == _information_T; // @[Lookup.scala 31:38]
  wire [31:0] _information_T_6 = io_in_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _information_T_7 = 32'h67 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_9 = 32'h63 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_11 = 32'h1063 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_13 = 32'h4063 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_15 = 32'h5063 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_17 = 32'h6063 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_19 = 32'h7063 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_21 = 32'h3 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_23 = 32'h1003 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_25 = 32'h2003 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_27 = 32'h4003 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_29 = 32'h5003 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_31 = 32'h23 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_33 = 32'h1023 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_35 = 32'h2023 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_37 = 32'h13 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_39 = 32'h2013 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_41 = 32'h3013 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_43 = 32'h4013 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_45 = 32'h6013 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_47 = 32'h7013 == _information_T_6; // @[Lookup.scala 31:38]
  wire [31:0] _information_T_48 = io_in_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _information_T_49 = 32'h1013 == _information_T_48; // @[Lookup.scala 31:38]
  wire  _information_T_51 = 32'h5013 == _information_T_48; // @[Lookup.scala 31:38]
  wire  _information_T_53 = 32'h40005013 == _information_T_48; // @[Lookup.scala 31:38]
  wire [31:0] _information_T_54 = io_in_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _information_T_55 = 32'h33 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_57 = 32'h40000033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_59 = 32'h1033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_61 = 32'h2033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_63 = 32'h3033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_65 = 32'h4033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_67 = 32'h5033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_69 = 32'h40005033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_71 = 32'h6033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_73 = 32'h7033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_75 = 32'h1b == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_77 = 32'h101b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_79 = 32'h501b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_81 = 32'h4000501b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_83 = 32'h3b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_85 = 32'h4000003b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_87 = 32'h103b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_89 = 32'h503b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_91 = 32'h4000503b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_93 = 32'h6003 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_95 = 32'h3003 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_97 = 32'h3023 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_99 = 32'h2000033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_101 = 32'h2001033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_103 = 32'h2002033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_105 = 32'h2003033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_107 = 32'h2004033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_109 = 32'h2005033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_111 = 32'h2006033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_113 = 32'h2007033 == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_115 = 32'h200003b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_117 = 32'h200403b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_119 = 32'h200503b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_121 = 32'h200603b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_123 = 32'h200703b == _information_T_54; // @[Lookup.scala 31:38]
  wire  _information_T_125 = 32'h100f == io_in_inst; // @[Lookup.scala 31:38]
  wire  _information_T_127 = 32'h1073 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_129 = 32'h2073 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_131 = 32'h3073 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_133 = 32'h5073 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_135 = 32'h6073 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_137 = 32'h7073 == _information_T_6; // @[Lookup.scala 31:38]
  wire  _information_T_139 = 32'h73 == io_in_inst; // @[Lookup.scala 31:38]
  wire  _information_T_141 = 32'h30200073 == io_in_inst; // @[Lookup.scala 31:38]
  wire [2:0] _information_T_221 = _information_T_139 ? 3'h1 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_222 = _information_T_137 ? 3'h1 : _information_T_221; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_223 = _information_T_135 ? 3'h1 : _information_T_222; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_224 = _information_T_133 ? 3'h1 : _information_T_223; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_225 = _information_T_131 ? 3'h1 : _information_T_224; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_226 = _information_T_129 ? 3'h1 : _information_T_225; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_227 = _information_T_127 ? 3'h1 : _information_T_226; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_228 = _information_T_125 ? 3'h1 : _information_T_227; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_229 = _information_T_123 ? 3'h0 : _information_T_228; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_230 = _information_T_121 ? 3'h0 : _information_T_229; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_231 = _information_T_119 ? 3'h0 : _information_T_230; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_232 = _information_T_117 ? 3'h0 : _information_T_231; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_233 = _information_T_115 ? 3'h0 : _information_T_232; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_234 = _information_T_113 ? 3'h0 : _information_T_233; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_235 = _information_T_111 ? 3'h0 : _information_T_234; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_236 = _information_T_109 ? 3'h0 : _information_T_235; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_237 = _information_T_107 ? 3'h0 : _information_T_236; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_238 = _information_T_105 ? 3'h0 : _information_T_237; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_239 = _information_T_103 ? 3'h0 : _information_T_238; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_240 = _information_T_101 ? 3'h0 : _information_T_239; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_241 = _information_T_99 ? 3'h0 : _information_T_240; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_242 = _information_T_97 ? 3'h2 : _information_T_241; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_243 = _information_T_95 ? 3'h1 : _information_T_242; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_244 = _information_T_93 ? 3'h1 : _information_T_243; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_245 = _information_T_91 ? 3'h0 : _information_T_244; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_246 = _information_T_89 ? 3'h0 : _information_T_245; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_247 = _information_T_87 ? 3'h0 : _information_T_246; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_248 = _information_T_85 ? 3'h0 : _information_T_247; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_249 = _information_T_83 ? 3'h0 : _information_T_248; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_250 = _information_T_81 ? 3'h1 : _information_T_249; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_251 = _information_T_79 ? 3'h1 : _information_T_250; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_252 = _information_T_77 ? 3'h1 : _information_T_251; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_253 = _information_T_75 ? 3'h1 : _information_T_252; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_254 = _information_T_73 ? 3'h0 : _information_T_253; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_255 = _information_T_71 ? 3'h0 : _information_T_254; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_256 = _information_T_69 ? 3'h0 : _information_T_255; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_257 = _information_T_67 ? 3'h0 : _information_T_256; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_258 = _information_T_65 ? 3'h0 : _information_T_257; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_259 = _information_T_63 ? 3'h0 : _information_T_258; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_260 = _information_T_61 ? 3'h0 : _information_T_259; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_261 = _information_T_59 ? 3'h0 : _information_T_260; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_262 = _information_T_57 ? 3'h0 : _information_T_261; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_263 = _information_T_55 ? 3'h0 : _information_T_262; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_264 = _information_T_53 ? 3'h1 : _information_T_263; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_265 = _information_T_51 ? 3'h1 : _information_T_264; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_266 = _information_T_49 ? 3'h1 : _information_T_265; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_267 = _information_T_47 ? 3'h1 : _information_T_266; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_268 = _information_T_45 ? 3'h1 : _information_T_267; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_269 = _information_T_43 ? 3'h1 : _information_T_268; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_270 = _information_T_41 ? 3'h1 : _information_T_269; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_271 = _information_T_39 ? 3'h1 : _information_T_270; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_272 = _information_T_37 ? 3'h1 : _information_T_271; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_273 = _information_T_35 ? 3'h2 : _information_T_272; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_274 = _information_T_33 ? 3'h2 : _information_T_273; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_275 = _information_T_31 ? 3'h2 : _information_T_274; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_276 = _information_T_29 ? 3'h1 : _information_T_275; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_277 = _information_T_27 ? 3'h1 : _information_T_276; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_278 = _information_T_25 ? 3'h1 : _information_T_277; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_279 = _information_T_23 ? 3'h1 : _information_T_278; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_280 = _information_T_21 ? 3'h1 : _information_T_279; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_281 = _information_T_19 ? 3'h3 : _information_T_280; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_282 = _information_T_17 ? 3'h3 : _information_T_281; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_283 = _information_T_15 ? 3'h3 : _information_T_282; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_284 = _information_T_13 ? 3'h3 : _information_T_283; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_285 = _information_T_11 ? 3'h3 : _information_T_284; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_286 = _information_T_9 ? 3'h3 : _information_T_285; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_287 = _information_T_7 ? 3'h1 : _information_T_286; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_288 = _information_T_5 ? 3'h5 : _information_T_287; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_289 = _information_T_3 ? 3'h4 : _information_T_288; // @[Lookup.scala 33:37]
  wire [2:0] information_1 = _information_T_1 ? 3'h4 : _information_T_289; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_292 = _information_T_141 ? 3'h3 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_293 = _information_T_139 ? 3'h3 : _information_T_292; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_294 = _information_T_137 ? 3'h3 : _information_T_293; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_295 = _information_T_135 ? 3'h3 : _information_T_294; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_296 = _information_T_133 ? 3'h3 : _information_T_295; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_297 = _information_T_131 ? 3'h3 : _information_T_296; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_298 = _information_T_129 ? 3'h3 : _information_T_297; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_299 = _information_T_127 ? 3'h3 : _information_T_298; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_300 = _information_T_125 ? 3'h3 : _information_T_299; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_301 = _information_T_123 ? 3'h4 : _information_T_300; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_302 = _information_T_121 ? 3'h4 : _information_T_301; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_303 = _information_T_119 ? 3'h4 : _information_T_302; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_304 = _information_T_117 ? 3'h4 : _information_T_303; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_305 = _information_T_115 ? 3'h4 : _information_T_304; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_306 = _information_T_113 ? 3'h4 : _information_T_305; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_307 = _information_T_111 ? 3'h4 : _information_T_306; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_308 = _information_T_109 ? 3'h4 : _information_T_307; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_309 = _information_T_107 ? 3'h4 : _information_T_308; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_310 = _information_T_105 ? 3'h4 : _information_T_309; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_311 = _information_T_103 ? 3'h4 : _information_T_310; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_312 = _information_T_101 ? 3'h4 : _information_T_311; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_313 = _information_T_99 ? 3'h4 : _information_T_312; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_314 = _information_T_97 ? 3'h2 : _information_T_313; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_315 = _information_T_95 ? 3'h2 : _information_T_314; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_316 = _information_T_93 ? 3'h2 : _information_T_315; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_317 = _information_T_91 ? 3'h0 : _information_T_316; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_318 = _information_T_89 ? 3'h0 : _information_T_317; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_319 = _information_T_87 ? 3'h0 : _information_T_318; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_320 = _information_T_85 ? 3'h0 : _information_T_319; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_321 = _information_T_83 ? 3'h0 : _information_T_320; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_322 = _information_T_81 ? 3'h0 : _information_T_321; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_323 = _information_T_79 ? 3'h0 : _information_T_322; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_324 = _information_T_77 ? 3'h0 : _information_T_323; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_325 = _information_T_75 ? 3'h0 : _information_T_324; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_326 = _information_T_73 ? 3'h0 : _information_T_325; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_327 = _information_T_71 ? 3'h0 : _information_T_326; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_328 = _information_T_69 ? 3'h0 : _information_T_327; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_329 = _information_T_67 ? 3'h0 : _information_T_328; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_330 = _information_T_65 ? 3'h0 : _information_T_329; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_331 = _information_T_63 ? 3'h0 : _information_T_330; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_332 = _information_T_61 ? 3'h0 : _information_T_331; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_333 = _information_T_59 ? 3'h0 : _information_T_332; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_334 = _information_T_57 ? 3'h0 : _information_T_333; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_335 = _information_T_55 ? 3'h0 : _information_T_334; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_336 = _information_T_53 ? 3'h0 : _information_T_335; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_337 = _information_T_51 ? 3'h0 : _information_T_336; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_338 = _information_T_49 ? 3'h0 : _information_T_337; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_339 = _information_T_47 ? 3'h0 : _information_T_338; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_340 = _information_T_45 ? 3'h0 : _information_T_339; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_341 = _information_T_43 ? 3'h0 : _information_T_340; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_342 = _information_T_41 ? 3'h0 : _information_T_341; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_343 = _information_T_39 ? 3'h0 : _information_T_342; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_344 = _information_T_37 ? 3'h0 : _information_T_343; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_345 = _information_T_35 ? 3'h2 : _information_T_344; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_346 = _information_T_33 ? 3'h2 : _information_T_345; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_347 = _information_T_31 ? 3'h2 : _information_T_346; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_348 = _information_T_29 ? 3'h2 : _information_T_347; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_349 = _information_T_27 ? 3'h2 : _information_T_348; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_350 = _information_T_25 ? 3'h2 : _information_T_349; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_351 = _information_T_23 ? 3'h2 : _information_T_350; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_352 = _information_T_21 ? 3'h2 : _information_T_351; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_353 = _information_T_19 ? 3'h1 : _information_T_352; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_354 = _information_T_17 ? 3'h1 : _information_T_353; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_355 = _information_T_15 ? 3'h1 : _information_T_354; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_356 = _information_T_13 ? 3'h1 : _information_T_355; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_357 = _information_T_11 ? 3'h1 : _information_T_356; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_358 = _information_T_9 ? 3'h1 : _information_T_357; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_359 = _information_T_7 ? 3'h1 : _information_T_358; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_360 = _information_T_5 ? 3'h1 : _information_T_359; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_361 = _information_T_3 ? 3'h0 : _information_T_360; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_389 = _information_T_91 ? 5'ha : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_390 = _information_T_89 ? 5'h9 : _information_T_389; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_391 = _information_T_87 ? 5'h8 : _information_T_390; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_392 = _information_T_85 ? 5'h2 : _information_T_391; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_393 = _information_T_83 ? 5'h1 : _information_T_392; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_394 = _information_T_81 ? 5'ha : _information_T_393; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_395 = _information_T_79 ? 5'h9 : _information_T_394; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_396 = _information_T_77 ? 5'h8 : _information_T_395; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_397 = _information_T_75 ? 5'h1 : _information_T_396; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_398 = _information_T_73 ? 5'h3 : _information_T_397; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_399 = _information_T_71 ? 5'h4 : _information_T_398; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_400 = _information_T_69 ? 5'ha : _information_T_399; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_401 = _information_T_67 ? 5'h9 : _information_T_400; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_402 = _information_T_65 ? 5'h5 : _information_T_401; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_403 = _information_T_63 ? 5'h7 : _information_T_402; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_404 = _information_T_61 ? 5'h6 : _information_T_403; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_405 = _information_T_59 ? 5'h8 : _information_T_404; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_406 = _information_T_57 ? 5'h2 : _information_T_405; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_407 = _information_T_55 ? 5'h1 : _information_T_406; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_408 = _information_T_53 ? 5'ha : _information_T_407; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_409 = _information_T_51 ? 5'h9 : _information_T_408; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_410 = _information_T_49 ? 5'h8 : _information_T_409; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_411 = _information_T_47 ? 5'h3 : _information_T_410; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_412 = _information_T_45 ? 5'h4 : _information_T_411; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_413 = _information_T_43 ? 5'h5 : _information_T_412; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_414 = _information_T_41 ? 5'h7 : _information_T_413; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_415 = _information_T_39 ? 5'h6 : _information_T_414; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_416 = _information_T_37 ? 5'h1 : _information_T_415; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_417 = _information_T_35 ? 5'h0 : _information_T_416; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_418 = _information_T_33 ? 5'h0 : _information_T_417; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_419 = _information_T_31 ? 5'h0 : _information_T_418; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_420 = _information_T_29 ? 5'h0 : _information_T_419; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_421 = _information_T_27 ? 5'h0 : _information_T_420; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_422 = _information_T_25 ? 5'h0 : _information_T_421; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_423 = _information_T_23 ? 5'h0 : _information_T_422; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_424 = _information_T_21 ? 5'h0 : _information_T_423; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_425 = _information_T_19 ? 5'h0 : _information_T_424; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_426 = _information_T_17 ? 5'h0 : _information_T_425; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_427 = _information_T_15 ? 5'h0 : _information_T_426; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_428 = _information_T_13 ? 5'h0 : _information_T_427; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_429 = _information_T_11 ? 5'h0 : _information_T_428; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_430 = _information_T_9 ? 5'h0 : _information_T_429; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_431 = _information_T_7 ? 5'h0 : _information_T_430; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_432 = _information_T_5 ? 5'h0 : _information_T_431; // @[Lookup.scala 33:37]
  wire [4:0] _information_T_433 = _information_T_3 ? 5'h1 : _information_T_432; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_497 = _information_T_19 ? 4'h8 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_498 = _information_T_17 ? 4'h7 : _information_T_497; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_499 = _information_T_15 ? 4'h6 : _information_T_498; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_500 = _information_T_13 ? 4'h5 : _information_T_499; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_501 = _information_T_11 ? 4'h4 : _information_T_500; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_502 = _information_T_9 ? 4'h3 : _information_T_501; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_503 = _information_T_7 ? 4'h2 : _information_T_502; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_504 = _information_T_5 ? 4'h1 : _information_T_503; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_505 = _information_T_3 ? 4'h0 : _information_T_504; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_530 = _information_T_97 ? 4'hb : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_531 = _information_T_95 ? 4'ha : _information_T_530; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_532 = _information_T_93 ? 4'h9 : _information_T_531; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_533 = _information_T_91 ? 4'h0 : _information_T_532; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_534 = _information_T_89 ? 4'h0 : _information_T_533; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_535 = _information_T_87 ? 4'h0 : _information_T_534; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_536 = _information_T_85 ? 4'h0 : _information_T_535; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_537 = _information_T_83 ? 4'h0 : _information_T_536; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_538 = _information_T_81 ? 4'h0 : _information_T_537; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_539 = _information_T_79 ? 4'h0 : _information_T_538; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_540 = _information_T_77 ? 4'h0 : _information_T_539; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_541 = _information_T_75 ? 4'h0 : _information_T_540; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_542 = _information_T_73 ? 4'h0 : _information_T_541; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_543 = _information_T_71 ? 4'h0 : _information_T_542; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_544 = _information_T_69 ? 4'h0 : _information_T_543; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_545 = _information_T_67 ? 4'h0 : _information_T_544; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_546 = _information_T_65 ? 4'h0 : _information_T_545; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_547 = _information_T_63 ? 4'h0 : _information_T_546; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_548 = _information_T_61 ? 4'h0 : _information_T_547; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_549 = _information_T_59 ? 4'h0 : _information_T_548; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_550 = _information_T_57 ? 4'h0 : _information_T_549; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_551 = _information_T_55 ? 4'h0 : _information_T_550; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_552 = _information_T_53 ? 4'h0 : _information_T_551; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_553 = _information_T_51 ? 4'h0 : _information_T_552; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_554 = _information_T_49 ? 4'h0 : _information_T_553; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_555 = _information_T_47 ? 4'h0 : _information_T_554; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_556 = _information_T_45 ? 4'h0 : _information_T_555; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_557 = _information_T_43 ? 4'h0 : _information_T_556; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_558 = _information_T_41 ? 4'h0 : _information_T_557; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_559 = _information_T_39 ? 4'h0 : _information_T_558; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_560 = _information_T_37 ? 4'h0 : _information_T_559; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_561 = _information_T_35 ? 4'h8 : _information_T_560; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_562 = _information_T_33 ? 4'h7 : _information_T_561; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_563 = _information_T_31 ? 4'h6 : _information_T_562; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_564 = _information_T_29 ? 4'h5 : _information_T_563; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_565 = _information_T_27 ? 4'h4 : _information_T_564; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_566 = _information_T_25 ? 4'h3 : _information_T_565; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_567 = _information_T_23 ? 4'h2 : _information_T_566; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_568 = _information_T_21 ? 4'h1 : _information_T_567; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_569 = _information_T_19 ? 4'h0 : _information_T_568; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_570 = _information_T_17 ? 4'h0 : _information_T_569; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_571 = _information_T_15 ? 4'h0 : _information_T_570; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_572 = _information_T_13 ? 4'h0 : _information_T_571; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_573 = _information_T_11 ? 4'h0 : _information_T_572; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_574 = _information_T_9 ? 4'h0 : _information_T_573; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_575 = _information_T_7 ? 4'h0 : _information_T_574; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_576 = _information_T_5 ? 4'h0 : _information_T_575; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_577 = _information_T_3 ? 4'h0 : _information_T_576; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_580 = _information_T_141 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_581 = _information_T_139 ? 3'h4 : _information_T_580; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_582 = _information_T_137 ? 3'h3 : _information_T_581; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_583 = _information_T_135 ? 3'h2 : _information_T_582; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_584 = _information_T_133 ? 3'h1 : _information_T_583; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_585 = _information_T_131 ? 3'h3 : _information_T_584; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_586 = _information_T_129 ? 3'h2 : _information_T_585; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_587 = _information_T_127 ? 3'h1 : _information_T_586; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_588 = _information_T_125 ? 3'h6 : _information_T_587; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_589 = _information_T_123 ? 3'h0 : _information_T_588; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_590 = _information_T_121 ? 3'h0 : _information_T_589; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_591 = _information_T_119 ? 3'h0 : _information_T_590; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_592 = _information_T_117 ? 3'h0 : _information_T_591; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_593 = _information_T_115 ? 3'h0 : _information_T_592; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_594 = _information_T_113 ? 3'h0 : _information_T_593; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_595 = _information_T_111 ? 3'h0 : _information_T_594; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_596 = _information_T_109 ? 3'h0 : _information_T_595; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_597 = _information_T_107 ? 3'h0 : _information_T_596; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_598 = _information_T_105 ? 3'h0 : _information_T_597; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_599 = _information_T_103 ? 3'h0 : _information_T_598; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_600 = _information_T_101 ? 3'h0 : _information_T_599; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_601 = _information_T_99 ? 3'h0 : _information_T_600; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_602 = _information_T_97 ? 3'h0 : _information_T_601; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_603 = _information_T_95 ? 3'h0 : _information_T_602; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_604 = _information_T_93 ? 3'h0 : _information_T_603; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_605 = _information_T_91 ? 3'h0 : _information_T_604; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_606 = _information_T_89 ? 3'h0 : _information_T_605; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_607 = _information_T_87 ? 3'h0 : _information_T_606; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_608 = _information_T_85 ? 3'h0 : _information_T_607; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_609 = _information_T_83 ? 3'h0 : _information_T_608; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_610 = _information_T_81 ? 3'h0 : _information_T_609; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_611 = _information_T_79 ? 3'h0 : _information_T_610; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_612 = _information_T_77 ? 3'h0 : _information_T_611; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_613 = _information_T_75 ? 3'h0 : _information_T_612; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_614 = _information_T_73 ? 3'h0 : _information_T_613; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_615 = _information_T_71 ? 3'h0 : _information_T_614; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_616 = _information_T_69 ? 3'h0 : _information_T_615; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_617 = _information_T_67 ? 3'h0 : _information_T_616; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_618 = _information_T_65 ? 3'h0 : _information_T_617; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_619 = _information_T_63 ? 3'h0 : _information_T_618; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_620 = _information_T_61 ? 3'h0 : _information_T_619; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_621 = _information_T_59 ? 3'h0 : _information_T_620; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_622 = _information_T_57 ? 3'h0 : _information_T_621; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_623 = _information_T_55 ? 3'h0 : _information_T_622; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_624 = _information_T_53 ? 3'h0 : _information_T_623; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_625 = _information_T_51 ? 3'h0 : _information_T_624; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_626 = _information_T_49 ? 3'h0 : _information_T_625; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_627 = _information_T_47 ? 3'h0 : _information_T_626; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_628 = _information_T_45 ? 3'h0 : _information_T_627; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_629 = _information_T_43 ? 3'h0 : _information_T_628; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_630 = _information_T_41 ? 3'h0 : _information_T_629; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_631 = _information_T_39 ? 3'h0 : _information_T_630; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_632 = _information_T_37 ? 3'h0 : _information_T_631; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_633 = _information_T_35 ? 3'h0 : _information_T_632; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_634 = _information_T_33 ? 3'h0 : _information_T_633; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_635 = _information_T_31 ? 3'h0 : _information_T_634; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_636 = _information_T_29 ? 3'h0 : _information_T_635; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_637 = _information_T_27 ? 3'h0 : _information_T_636; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_638 = _information_T_25 ? 3'h0 : _information_T_637; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_639 = _information_T_23 ? 3'h0 : _information_T_638; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_640 = _information_T_21 ? 3'h0 : _information_T_639; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_641 = _information_T_19 ? 3'h0 : _information_T_640; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_642 = _information_T_17 ? 3'h0 : _information_T_641; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_643 = _information_T_15 ? 3'h0 : _information_T_642; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_644 = _information_T_13 ? 3'h0 : _information_T_643; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_645 = _information_T_11 ? 3'h0 : _information_T_644; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_646 = _information_T_9 ? 3'h0 : _information_T_645; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_647 = _information_T_7 ? 3'h0 : _information_T_646; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_648 = _information_T_5 ? 3'h0 : _information_T_647; // @[Lookup.scala 33:37]
  wire [2:0] _information_T_649 = _information_T_3 ? 3'h0 : _information_T_648; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_661 = _information_T_123 ? 4'h8 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_662 = _information_T_121 ? 4'h7 : _information_T_661; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_663 = _information_T_119 ? 4'h6 : _information_T_662; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_664 = _information_T_117 ? 4'h5 : _information_T_663; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_665 = _information_T_115 ? 4'h1 : _information_T_664; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_666 = _information_T_113 ? 4'h8 : _information_T_665; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_667 = _information_T_111 ? 4'h7 : _information_T_666; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_668 = _information_T_109 ? 4'h6 : _information_T_667; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_669 = _information_T_107 ? 4'h5 : _information_T_668; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_670 = _information_T_105 ? 4'h4 : _information_T_669; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_671 = _information_T_103 ? 4'h3 : _information_T_670; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_672 = _information_T_101 ? 4'h2 : _information_T_671; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_673 = _information_T_99 ? 4'h1 : _information_T_672; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_674 = _information_T_97 ? 4'h0 : _information_T_673; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_675 = _information_T_95 ? 4'h0 : _information_T_674; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_676 = _information_T_93 ? 4'h0 : _information_T_675; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_677 = _information_T_91 ? 4'h0 : _information_T_676; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_678 = _information_T_89 ? 4'h0 : _information_T_677; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_679 = _information_T_87 ? 4'h0 : _information_T_678; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_680 = _information_T_85 ? 4'h0 : _information_T_679; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_681 = _information_T_83 ? 4'h0 : _information_T_680; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_682 = _information_T_81 ? 4'h0 : _information_T_681; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_683 = _information_T_79 ? 4'h0 : _information_T_682; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_684 = _information_T_77 ? 4'h0 : _information_T_683; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_685 = _information_T_75 ? 4'h0 : _information_T_684; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_686 = _information_T_73 ? 4'h0 : _information_T_685; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_687 = _information_T_71 ? 4'h0 : _information_T_686; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_688 = _information_T_69 ? 4'h0 : _information_T_687; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_689 = _information_T_67 ? 4'h0 : _information_T_688; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_690 = _information_T_65 ? 4'h0 : _information_T_689; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_691 = _information_T_63 ? 4'h0 : _information_T_690; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_692 = _information_T_61 ? 4'h0 : _information_T_691; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_693 = _information_T_59 ? 4'h0 : _information_T_692; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_694 = _information_T_57 ? 4'h0 : _information_T_693; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_695 = _information_T_55 ? 4'h0 : _information_T_694; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_696 = _information_T_53 ? 4'h0 : _information_T_695; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_697 = _information_T_51 ? 4'h0 : _information_T_696; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_698 = _information_T_49 ? 4'h0 : _information_T_697; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_699 = _information_T_47 ? 4'h0 : _information_T_698; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_700 = _information_T_45 ? 4'h0 : _information_T_699; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_701 = _information_T_43 ? 4'h0 : _information_T_700; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_702 = _information_T_41 ? 4'h0 : _information_T_701; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_703 = _information_T_39 ? 4'h0 : _information_T_702; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_704 = _information_T_37 ? 4'h0 : _information_T_703; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_705 = _information_T_35 ? 4'h0 : _information_T_704; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_706 = _information_T_33 ? 4'h0 : _information_T_705; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_707 = _information_T_31 ? 4'h0 : _information_T_706; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_708 = _information_T_29 ? 4'h0 : _information_T_707; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_709 = _information_T_27 ? 4'h0 : _information_T_708; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_710 = _information_T_25 ? 4'h0 : _information_T_709; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_711 = _information_T_23 ? 4'h0 : _information_T_710; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_712 = _information_T_21 ? 4'h0 : _information_T_711; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_713 = _information_T_19 ? 4'h0 : _information_T_712; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_714 = _information_T_17 ? 4'h0 : _information_T_713; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_715 = _information_T_15 ? 4'h0 : _information_T_714; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_716 = _information_T_13 ? 4'h0 : _information_T_715; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_717 = _information_T_11 ? 4'h0 : _information_T_716; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_718 = _information_T_9 ? 4'h0 : _information_T_717; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_719 = _information_T_7 ? 4'h0 : _information_T_718; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_720 = _information_T_5 ? 4'h0 : _information_T_719; // @[Lookup.scala 33:37]
  wire [3:0] _information_T_721 = _information_T_3 ? 4'h0 : _information_T_720; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_726 = _information_T_137 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_727 = _information_T_135 ? 2'h3 : _information_T_726; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_728 = _information_T_133 ? 2'h3 : _information_T_727; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_729 = _information_T_131 ? 2'h2 : _information_T_728; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_730 = _information_T_129 ? 2'h2 : _information_T_729; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_731 = _information_T_127 ? 2'h2 : _information_T_730; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_732 = _information_T_125 ? 2'h0 : _information_T_731; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_733 = _information_T_123 ? 2'h2 : _information_T_732; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_734 = _information_T_121 ? 2'h2 : _information_T_733; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_735 = _information_T_119 ? 2'h2 : _information_T_734; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_736 = _information_T_117 ? 2'h2 : _information_T_735; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_737 = _information_T_115 ? 2'h2 : _information_T_736; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_738 = _information_T_113 ? 2'h2 : _information_T_737; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_739 = _information_T_111 ? 2'h2 : _information_T_738; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_740 = _information_T_109 ? 2'h2 : _information_T_739; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_741 = _information_T_107 ? 2'h2 : _information_T_740; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_742 = _information_T_105 ? 2'h2 : _information_T_741; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_743 = _information_T_103 ? 2'h2 : _information_T_742; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_744 = _information_T_101 ? 2'h2 : _information_T_743; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_745 = _information_T_99 ? 2'h2 : _information_T_744; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_746 = _information_T_97 ? 2'h2 : _information_T_745; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_747 = _information_T_95 ? 2'h2 : _information_T_746; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_748 = _information_T_93 ? 2'h2 : _information_T_747; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_749 = _information_T_91 ? 2'h2 : _information_T_748; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_750 = _information_T_89 ? 2'h2 : _information_T_749; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_751 = _information_T_87 ? 2'h2 : _information_T_750; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_752 = _information_T_85 ? 2'h2 : _information_T_751; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_753 = _information_T_83 ? 2'h2 : _information_T_752; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_754 = _information_T_81 ? 2'h2 : _information_T_753; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_755 = _information_T_79 ? 2'h2 : _information_T_754; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_756 = _information_T_77 ? 2'h2 : _information_T_755; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_757 = _information_T_75 ? 2'h2 : _information_T_756; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_758 = _information_T_73 ? 2'h2 : _information_T_757; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_759 = _information_T_71 ? 2'h2 : _information_T_758; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_760 = _information_T_69 ? 2'h2 : _information_T_759; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_761 = _information_T_67 ? 2'h2 : _information_T_760; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_762 = _information_T_65 ? 2'h2 : _information_T_761; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_763 = _information_T_63 ? 2'h2 : _information_T_762; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_764 = _information_T_61 ? 2'h2 : _information_T_763; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_765 = _information_T_59 ? 2'h2 : _information_T_764; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_766 = _information_T_57 ? 2'h2 : _information_T_765; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_767 = _information_T_55 ? 2'h2 : _information_T_766; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_768 = _information_T_53 ? 2'h2 : _information_T_767; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_769 = _information_T_51 ? 2'h2 : _information_T_768; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_770 = _information_T_49 ? 2'h2 : _information_T_769; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_771 = _information_T_47 ? 2'h2 : _information_T_770; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_772 = _information_T_45 ? 2'h2 : _information_T_771; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_773 = _information_T_43 ? 2'h2 : _information_T_772; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_774 = _information_T_41 ? 2'h2 : _information_T_773; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_775 = _information_T_39 ? 2'h2 : _information_T_774; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_776 = _information_T_37 ? 2'h2 : _information_T_775; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_777 = _information_T_35 ? 2'h2 : _information_T_776; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_778 = _information_T_33 ? 2'h2 : _information_T_777; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_779 = _information_T_31 ? 2'h2 : _information_T_778; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_780 = _information_T_29 ? 2'h2 : _information_T_779; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_781 = _information_T_27 ? 2'h2 : _information_T_780; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_782 = _information_T_25 ? 2'h2 : _information_T_781; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_783 = _information_T_23 ? 2'h2 : _information_T_782; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_784 = _information_T_21 ? 2'h2 : _information_T_783; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_785 = _information_T_19 ? 2'h2 : _information_T_784; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_786 = _information_T_17 ? 2'h2 : _information_T_785; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_787 = _information_T_15 ? 2'h2 : _information_T_786; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_788 = _information_T_13 ? 2'h2 : _information_T_787; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_789 = _information_T_11 ? 2'h2 : _information_T_788; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_790 = _information_T_9 ? 2'h2 : _information_T_789; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_791 = _information_T_7 ? 2'h2 : _information_T_790; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_792 = _information_T_5 ? 2'h1 : _information_T_791; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_793 = _information_T_3 ? 2'h1 : _information_T_792; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_805 = _information_T_123 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_806 = _information_T_121 ? 2'h2 : _information_T_805; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_807 = _information_T_119 ? 2'h2 : _information_T_806; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_808 = _information_T_117 ? 2'h2 : _information_T_807; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_809 = _information_T_115 ? 2'h2 : _information_T_808; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_810 = _information_T_113 ? 2'h2 : _information_T_809; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_811 = _information_T_111 ? 2'h2 : _information_T_810; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_812 = _information_T_109 ? 2'h2 : _information_T_811; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_813 = _information_T_107 ? 2'h2 : _information_T_812; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_814 = _information_T_105 ? 2'h2 : _information_T_813; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_815 = _information_T_103 ? 2'h2 : _information_T_814; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_816 = _information_T_101 ? 2'h2 : _information_T_815; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_817 = _information_T_99 ? 2'h2 : _information_T_816; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_818 = _information_T_97 ? 2'h3 : _information_T_817; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_819 = _information_T_95 ? 2'h3 : _information_T_818; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_820 = _information_T_93 ? 2'h3 : _information_T_819; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_821 = _information_T_91 ? 2'h2 : _information_T_820; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_822 = _information_T_89 ? 2'h2 : _information_T_821; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_823 = _information_T_87 ? 2'h2 : _information_T_822; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_824 = _information_T_85 ? 2'h2 : _information_T_823; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_825 = _information_T_83 ? 2'h2 : _information_T_824; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_826 = _information_T_81 ? 2'h3 : _information_T_825; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_827 = _information_T_79 ? 2'h3 : _information_T_826; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_828 = _information_T_77 ? 2'h3 : _information_T_827; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_829 = _information_T_75 ? 2'h3 : _information_T_828; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_830 = _information_T_73 ? 2'h2 : _information_T_829; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_831 = _information_T_71 ? 2'h2 : _information_T_830; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_832 = _information_T_69 ? 2'h2 : _information_T_831; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_833 = _information_T_67 ? 2'h2 : _information_T_832; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_834 = _information_T_65 ? 2'h2 : _information_T_833; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_835 = _information_T_63 ? 2'h2 : _information_T_834; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_836 = _information_T_61 ? 2'h2 : _information_T_835; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_837 = _information_T_59 ? 2'h2 : _information_T_836; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_838 = _information_T_57 ? 2'h2 : _information_T_837; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_839 = _information_T_55 ? 2'h2 : _information_T_838; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_840 = _information_T_53 ? 2'h3 : _information_T_839; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_841 = _information_T_51 ? 2'h3 : _information_T_840; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_842 = _information_T_49 ? 2'h3 : _information_T_841; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_843 = _information_T_47 ? 2'h3 : _information_T_842; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_844 = _information_T_45 ? 2'h3 : _information_T_843; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_845 = _information_T_43 ? 2'h3 : _information_T_844; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_846 = _information_T_41 ? 2'h3 : _information_T_845; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_847 = _information_T_39 ? 2'h3 : _information_T_846; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_848 = _information_T_37 ? 2'h3 : _information_T_847; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_849 = _information_T_35 ? 2'h3 : _information_T_848; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_850 = _information_T_33 ? 2'h3 : _information_T_849; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_851 = _information_T_31 ? 2'h3 : _information_T_850; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_852 = _information_T_29 ? 2'h3 : _information_T_851; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_853 = _information_T_27 ? 2'h3 : _information_T_852; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_854 = _information_T_25 ? 2'h3 : _information_T_853; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_855 = _information_T_23 ? 2'h3 : _information_T_854; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_856 = _information_T_21 ? 2'h3 : _information_T_855; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_857 = _information_T_19 ? 2'h2 : _information_T_856; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_858 = _information_T_17 ? 2'h2 : _information_T_857; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_859 = _information_T_15 ? 2'h2 : _information_T_858; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_860 = _information_T_13 ? 2'h2 : _information_T_859; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_861 = _information_T_11 ? 2'h2 : _information_T_860; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_862 = _information_T_9 ? 2'h2 : _information_T_861; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_863 = _information_T_7 ? 2'h3 : _information_T_862; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_864 = _information_T_5 ? 2'h3 : _information_T_863; // @[Lookup.scala 33:37]
  wire [1:0] _information_T_865 = _information_T_3 ? 2'h3 : _information_T_864; // @[Lookup.scala 33:37]
  wire  _information_T_876 = _information_T_125 ? 1'h0 : _information_T_127 | (_information_T_129 | (_information_T_131
     | (_information_T_133 | (_information_T_135 | _information_T_137)))); // @[Lookup.scala 33:37]
  wire  _information_T_890 = _information_T_97 ? 1'h0 : _information_T_99 | (_information_T_101 | (_information_T_103 |
    (_information_T_105 | (_information_T_107 | (_information_T_109 | (_information_T_111 | (_information_T_113 | (
    _information_T_115 | (_information_T_117 | (_information_T_119 | (_information_T_121 | (_information_T_123 |
    _information_T_876)))))))))))); // @[Lookup.scala 33:37]
  wire  _information_T_920 = _information_T_37 | (_information_T_39 | (_information_T_41 | (_information_T_43 | (
    _information_T_45 | (_information_T_47 | (_information_T_49 | (_information_T_51 | (_information_T_53 | (
    _information_T_55 | (_information_T_57 | (_information_T_59 | (_information_T_61 | (_information_T_63 | (
    _information_T_65 | (_information_T_67 | (_information_T_69 | (_information_T_71 | (_information_T_73 | (
    _information_T_75 | (_information_T_77 | (_information_T_79 | (_information_T_81 | (_information_T_83 | (
    _information_T_85 | (_information_T_87 | (_information_T_89 | (_information_T_91 | (_information_T_93 | (
    _information_T_95 | _information_T_890))))))))))))))))))))))))))))); // @[Lookup.scala 33:37]
  wire  _information_T_921 = _information_T_35 ? 1'h0 : _information_T_920; // @[Lookup.scala 33:37]
  wire  _information_T_922 = _information_T_33 ? 1'h0 : _information_T_921; // @[Lookup.scala 33:37]
  wire  _information_T_923 = _information_T_31 ? 1'h0 : _information_T_922; // @[Lookup.scala 33:37]
  wire  _information_T_929 = _information_T_19 ? 1'h0 : _information_T_21 | (_information_T_23 | (_information_T_25 | (
    _information_T_27 | (_information_T_29 | _information_T_923)))); // @[Lookup.scala 33:37]
  wire  _information_T_930 = _information_T_17 ? 1'h0 : _information_T_929; // @[Lookup.scala 33:37]
  wire  _information_T_931 = _information_T_15 ? 1'h0 : _information_T_930; // @[Lookup.scala 33:37]
  wire  _information_T_932 = _information_T_13 ? 1'h0 : _information_T_931; // @[Lookup.scala 33:37]
  wire  _information_T_933 = _information_T_11 ? 1'h0 : _information_T_932; // @[Lookup.scala 33:37]
  wire  _information_T_934 = _information_T_9 ? 1'h0 : _information_T_933; // @[Lookup.scala 33:37]
  wire  _information_T_954 = _information_T_113 ? 1'h0 : _information_T_115 | (_information_T_117 | (_information_T_119
     | (_information_T_121 | _information_T_123))); // @[Lookup.scala 33:37]
  wire  _information_T_955 = _information_T_111 ? 1'h0 : _information_T_954; // @[Lookup.scala 33:37]
  wire  _information_T_956 = _information_T_109 ? 1'h0 : _information_T_955; // @[Lookup.scala 33:37]
  wire  _information_T_957 = _information_T_107 ? 1'h0 : _information_T_956; // @[Lookup.scala 33:37]
  wire  _information_T_958 = _information_T_105 ? 1'h0 : _information_T_957; // @[Lookup.scala 33:37]
  wire  _information_T_959 = _information_T_103 ? 1'h0 : _information_T_958; // @[Lookup.scala 33:37]
  wire  _information_T_960 = _information_T_101 ? 1'h0 : _information_T_959; // @[Lookup.scala 33:37]
  wire  _information_T_961 = _information_T_99 ? 1'h0 : _information_T_960; // @[Lookup.scala 33:37]
  wire  _information_T_962 = _information_T_97 ? 1'h0 : _information_T_961; // @[Lookup.scala 33:37]
  wire  _information_T_963 = _information_T_95 ? 1'h0 : _information_T_962; // @[Lookup.scala 33:37]
  wire  _information_T_964 = _information_T_93 ? 1'h0 : _information_T_963; // @[Lookup.scala 33:37]
  wire  _information_T_974 = _information_T_73 ? 1'h0 : _information_T_75 | (_information_T_77 | (_information_T_79 | (
    _information_T_81 | (_information_T_83 | (_information_T_85 | (_information_T_87 | (_information_T_89 | (
    _information_T_91 | _information_T_964)))))))); // @[Lookup.scala 33:37]
  wire  _information_T_975 = _information_T_71 ? 1'h0 : _information_T_974; // @[Lookup.scala 33:37]
  wire  _information_T_976 = _information_T_69 ? 1'h0 : _information_T_975; // @[Lookup.scala 33:37]
  wire  _information_T_977 = _information_T_67 ? 1'h0 : _information_T_976; // @[Lookup.scala 33:37]
  wire  _information_T_978 = _information_T_65 ? 1'h0 : _information_T_977; // @[Lookup.scala 33:37]
  wire  _information_T_979 = _information_T_63 ? 1'h0 : _information_T_978; // @[Lookup.scala 33:37]
  wire  _information_T_980 = _information_T_61 ? 1'h0 : _information_T_979; // @[Lookup.scala 33:37]
  wire  _information_T_981 = _information_T_59 ? 1'h0 : _information_T_980; // @[Lookup.scala 33:37]
  wire  _information_T_982 = _information_T_57 ? 1'h0 : _information_T_981; // @[Lookup.scala 33:37]
  wire  _information_T_983 = _information_T_55 ? 1'h0 : _information_T_982; // @[Lookup.scala 33:37]
  wire  _information_T_984 = _information_T_53 ? 1'h0 : _information_T_983; // @[Lookup.scala 33:37]
  wire  _information_T_985 = _information_T_51 ? 1'h0 : _information_T_984; // @[Lookup.scala 33:37]
  wire  _information_T_986 = _information_T_49 ? 1'h0 : _information_T_985; // @[Lookup.scala 33:37]
  wire  _information_T_987 = _information_T_47 ? 1'h0 : _information_T_986; // @[Lookup.scala 33:37]
  wire  _information_T_988 = _information_T_45 ? 1'h0 : _information_T_987; // @[Lookup.scala 33:37]
  wire  _information_T_989 = _information_T_43 ? 1'h0 : _information_T_988; // @[Lookup.scala 33:37]
  wire  _information_T_990 = _information_T_41 ? 1'h0 : _information_T_989; // @[Lookup.scala 33:37]
  wire  _information_T_991 = _information_T_39 ? 1'h0 : _information_T_990; // @[Lookup.scala 33:37]
  wire  _information_T_992 = _information_T_37 ? 1'h0 : _information_T_991; // @[Lookup.scala 33:37]
  wire  _information_T_993 = _information_T_35 ? 1'h0 : _information_T_992; // @[Lookup.scala 33:37]
  wire  _information_T_994 = _information_T_33 ? 1'h0 : _information_T_993; // @[Lookup.scala 33:37]
  wire  _information_T_995 = _information_T_31 ? 1'h0 : _information_T_994; // @[Lookup.scala 33:37]
  wire  _information_T_996 = _information_T_29 ? 1'h0 : _information_T_995; // @[Lookup.scala 33:37]
  wire  _information_T_997 = _information_T_27 ? 1'h0 : _information_T_996; // @[Lookup.scala 33:37]
  wire  _information_T_998 = _information_T_25 ? 1'h0 : _information_T_997; // @[Lookup.scala 33:37]
  wire  _information_T_999 = _information_T_23 ? 1'h0 : _information_T_998; // @[Lookup.scala 33:37]
  wire  _information_T_1000 = _information_T_21 ? 1'h0 : _information_T_999; // @[Lookup.scala 33:37]
  wire  _information_T_1001 = _information_T_19 ? 1'h0 : _information_T_1000; // @[Lookup.scala 33:37]
  wire  _information_T_1002 = _information_T_17 ? 1'h0 : _information_T_1001; // @[Lookup.scala 33:37]
  wire  _information_T_1003 = _information_T_15 ? 1'h0 : _information_T_1002; // @[Lookup.scala 33:37]
  wire  _information_T_1004 = _information_T_13 ? 1'h0 : _information_T_1003; // @[Lookup.scala 33:37]
  wire  _information_T_1005 = _information_T_11 ? 1'h0 : _information_T_1004; // @[Lookup.scala 33:37]
  wire  _information_T_1006 = _information_T_9 ? 1'h0 : _information_T_1005; // @[Lookup.scala 33:37]
  wire  _information_T_1007 = _information_T_7 ? 1'h0 : _information_T_1006; // @[Lookup.scala 33:37]
  wire  _information_T_1008 = _information_T_5 ? 1'h0 : _information_T_1007; // @[Lookup.scala 33:37]
  wire  _information_T_1009 = _information_T_3 ? 1'h0 : _information_T_1008; // @[Lookup.scala 33:37]
  wire [63:0] _imm_T_1 = 3'h1 == information_1 ? imm_i : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_3 = 3'h2 == information_1 ? imm_s : _imm_T_1; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_5 = 3'h3 == information_1 ? imm_b : _imm_T_3; // @[Mux.scala 80:57]
  wire [63:0] _imm_T_7 = 3'h4 == information_1 ? imm_u : _imm_T_5; // @[Mux.scala 80:57]
  assign io_out_valid = io_in_valid; // @[IDU.scala 133:13]
  assign io_out_pc = io_in_pc; // @[IDU.scala 134:10]
  assign io_out_inst = io_in_inst; // @[IDU.scala 135:12]
  assign io_out_src1 = _information_T_1 ? 2'h0 : _information_T_793; // @[Lookup.scala 33:37]
  assign io_out_src2 = _information_T_1 ? 2'h3 : _information_T_865; // @[Lookup.scala 33:37]
  assign io_out_rs1 = io_in_inst[19:15]; // @[IDU.scala 121:14]
  assign io_out_rs2 = io_in_inst[24:20]; // @[IDU.scala 122:14]
  assign io_out_dest = io_in_inst[11:7]; // @[IDU.scala 123:15]
  assign io_out_imm = 3'h5 == information_1 ? imm_j : _imm_T_7; // @[Mux.scala 80:57]
  assign io_out_fu_type = _information_T_1 ? 3'h0 : _information_T_361; // @[Lookup.scala 33:37]
  assign io_out_bru_op = _information_T_1 ? 4'h0 : _information_T_505; // @[Lookup.scala 33:37]
  assign io_out_alu_op = _information_T_1 ? 5'h1 : _information_T_433; // @[Lookup.scala 33:37]
  assign io_out_lsu_op = _information_T_1 ? 4'h0 : _information_T_577; // @[Lookup.scala 33:37]
  assign io_out_csr_op = _information_T_1 ? 3'h0 : _information_T_649; // @[Lookup.scala 33:37]
  assign io_out_mdu_op = _information_T_1 ? 4'h0 : _information_T_721; // @[Lookup.scala 33:37]
  assign io_out_wen = _information_T_1 | (_information_T_3 | (_information_T_5 | (_information_T_7 | _information_T_934)
    )); // @[Lookup.scala 33:37]
  assign io_out_rv64 = _information_T_1 ? 1'h0 : _information_T_1009; // @[Lookup.scala 33:37]
  assign io_out_bp_br_taken = io_in_bp_br_taken; // @[IDU.scala 150:19]
  assign io_out_bp_br_target = io_in_bp_br_target; // @[IDU.scala 151:20]
  assign io_out_bp_br_type = io_in_bp_br_type; // @[IDU.scala 152:18]
endmodule
module IDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_0_valid,
  input  [31:0] io_in_bits_0_pc,
  input  [31:0] io_in_bits_0_inst,
  input         io_in_bits_0_bp_br_taken,
  input  [31:0] io_in_bits_0_bp_br_target,
  input  [1:0]  io_in_bits_0_bp_br_type,
  input         io_in_bits_1_valid,
  input  [31:0] io_in_bits_1_pc,
  input  [31:0] io_in_bits_1_inst,
  input         io_in_bits_1_bp_br_taken,
  input  [31:0] io_in_bits_1_bp_br_target,
  input  [1:0]  io_in_bits_1_bp_br_type,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_0_valid,
  output [31:0] io_out_bits_0_pc,
  output [31:0] io_out_bits_0_inst,
  output [1:0]  io_out_bits_0_src1,
  output [1:0]  io_out_bits_0_src2,
  output [4:0]  io_out_bits_0_rs1,
  output [4:0]  io_out_bits_0_rs2,
  output [4:0]  io_out_bits_0_dest,
  output [63:0] io_out_bits_0_imm,
  output [2:0]  io_out_bits_0_fu_type,
  output [3:0]  io_out_bits_0_bru_op,
  output [4:0]  io_out_bits_0_alu_op,
  output [3:0]  io_out_bits_0_lsu_op,
  output [2:0]  io_out_bits_0_csr_op,
  output [3:0]  io_out_bits_0_mdu_op,
  output        io_out_bits_0_wen,
  output        io_out_bits_0_rv64,
  output        io_out_bits_0_bp_br_taken,
  output [31:0] io_out_bits_0_bp_br_target,
  output [1:0]  io_out_bits_0_bp_br_type,
  output        io_out_bits_1_valid,
  output [31:0] io_out_bits_1_pc,
  output [31:0] io_out_bits_1_inst,
  output [1:0]  io_out_bits_1_src1,
  output [1:0]  io_out_bits_1_src2,
  output [4:0]  io_out_bits_1_rs1,
  output [4:0]  io_out_bits_1_rs2,
  output [4:0]  io_out_bits_1_dest,
  output [63:0] io_out_bits_1_imm,
  output [2:0]  io_out_bits_1_fu_type,
  output [3:0]  io_out_bits_1_bru_op,
  output [4:0]  io_out_bits_1_alu_op,
  output [3:0]  io_out_bits_1_lsu_op,
  output [2:0]  io_out_bits_1_csr_op,
  output [3:0]  io_out_bits_1_mdu_op,
  output        io_out_bits_1_wen,
  output        io_out_bits_1_rv64,
  output        io_out_bits_1_bp_br_taken,
  output [31:0] io_out_bits_1_bp_br_target,
  output [1:0]  io_out_bits_1_bp_br_type,
  input         frontend_reflush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  decode_entry_0_io_in_valid; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_0_io_in_pc; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_0_io_in_inst; // @[IDU.scala 163:30]
  wire  decode_entry_0_io_in_bp_br_taken; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_0_io_in_bp_br_target; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_0_io_in_bp_br_type; // @[IDU.scala 163:30]
  wire  decode_entry_0_io_out_valid; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_0_io_out_pc; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_0_io_out_inst; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_0_io_out_src1; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_0_io_out_src2; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_0_io_out_rs1; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_0_io_out_rs2; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_0_io_out_dest; // @[IDU.scala 163:30]
  wire [63:0] decode_entry_0_io_out_imm; // @[IDU.scala 163:30]
  wire [2:0] decode_entry_0_io_out_fu_type; // @[IDU.scala 163:30]
  wire [3:0] decode_entry_0_io_out_bru_op; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_0_io_out_alu_op; // @[IDU.scala 163:30]
  wire [3:0] decode_entry_0_io_out_lsu_op; // @[IDU.scala 163:30]
  wire [2:0] decode_entry_0_io_out_csr_op; // @[IDU.scala 163:30]
  wire [3:0] decode_entry_0_io_out_mdu_op; // @[IDU.scala 163:30]
  wire  decode_entry_0_io_out_wen; // @[IDU.scala 163:30]
  wire  decode_entry_0_io_out_rv64; // @[IDU.scala 163:30]
  wire  decode_entry_0_io_out_bp_br_taken; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_0_io_out_bp_br_target; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_0_io_out_bp_br_type; // @[IDU.scala 163:30]
  wire  decode_entry_1_io_in_valid; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_1_io_in_pc; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_1_io_in_inst; // @[IDU.scala 163:30]
  wire  decode_entry_1_io_in_bp_br_taken; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_1_io_in_bp_br_target; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_1_io_in_bp_br_type; // @[IDU.scala 163:30]
  wire  decode_entry_1_io_out_valid; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_1_io_out_pc; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_1_io_out_inst; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_1_io_out_src1; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_1_io_out_src2; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_1_io_out_rs1; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_1_io_out_rs2; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_1_io_out_dest; // @[IDU.scala 163:30]
  wire [63:0] decode_entry_1_io_out_imm; // @[IDU.scala 163:30]
  wire [2:0] decode_entry_1_io_out_fu_type; // @[IDU.scala 163:30]
  wire [3:0] decode_entry_1_io_out_bru_op; // @[IDU.scala 163:30]
  wire [4:0] decode_entry_1_io_out_alu_op; // @[IDU.scala 163:30]
  wire [3:0] decode_entry_1_io_out_lsu_op; // @[IDU.scala 163:30]
  wire [2:0] decode_entry_1_io_out_csr_op; // @[IDU.scala 163:30]
  wire [3:0] decode_entry_1_io_out_mdu_op; // @[IDU.scala 163:30]
  wire  decode_entry_1_io_out_wen; // @[IDU.scala 163:30]
  wire  decode_entry_1_io_out_rv64; // @[IDU.scala 163:30]
  wire  decode_entry_1_io_out_bp_br_taken; // @[IDU.scala 163:30]
  wire [31:0] decode_entry_1_io_out_bp_br_target; // @[IDU.scala 163:30]
  wire [1:0] decode_entry_1_io_out_bp_br_type; // @[IDU.scala 163:30]
  reg  conflict_decode_entry_valid; // @[IDU.scala 172:38]
  reg [31:0] conflict_decode_entry_pc; // @[IDU.scala 172:38]
  reg [31:0] conflict_decode_entry_inst; // @[IDU.scala 172:38]
  reg [1:0] conflict_decode_entry_src1; // @[IDU.scala 172:38]
  reg [1:0] conflict_decode_entry_src2; // @[IDU.scala 172:38]
  reg [4:0] conflict_decode_entry_rs1; // @[IDU.scala 172:38]
  reg [4:0] conflict_decode_entry_rs2; // @[IDU.scala 172:38]
  reg [4:0] conflict_decode_entry_dest; // @[IDU.scala 172:38]
  reg [63:0] conflict_decode_entry_imm; // @[IDU.scala 172:38]
  reg [2:0] conflict_decode_entry_fu_type; // @[IDU.scala 172:38]
  reg [3:0] conflict_decode_entry_bru_op; // @[IDU.scala 172:38]
  reg [4:0] conflict_decode_entry_alu_op; // @[IDU.scala 172:38]
  reg [3:0] conflict_decode_entry_lsu_op; // @[IDU.scala 172:38]
  reg [2:0] conflict_decode_entry_csr_op; // @[IDU.scala 172:38]
  reg [3:0] conflict_decode_entry_mdu_op; // @[IDU.scala 172:38]
  reg  conflict_decode_entry_wen; // @[IDU.scala 172:38]
  reg  conflict_decode_entry_rv64; // @[IDU.scala 172:38]
  reg  conflict_decode_entry_bp_br_taken; // @[IDU.scala 172:38]
  reg [31:0] conflict_decode_entry_bp_br_target; // @[IDU.scala 172:38]
  reg [1:0] conflict_decode_entry_bp_br_type; // @[IDU.scala 172:38]
  reg  had_conflict; // @[IDU.scala 174:29]
  wire  _self_reg_conflict_T_1 = decode_entry_1_io_out_rs1 != 5'h0; // @[IDU.scala 180:32]
  wire  _self_reg_conflict_T_2 = decode_entry_1_io_out_src1 == 2'h2 & _self_reg_conflict_T_1; // @[IDU.scala 179:64]
  wire  _self_reg_conflict_T_3 = decode_entry_1_io_out_rs1 == decode_entry_0_io_out_dest; // @[IDU.scala 181:32]
  wire  _self_reg_conflict_T_4 = _self_reg_conflict_T_2 & _self_reg_conflict_T_3; // @[IDU.scala 180:40]
  wire  _self_reg_conflict_T_5 = _self_reg_conflict_T_4 & decode_entry_0_io_out_wen; // @[IDU.scala 181:64]
  wire  _self_reg_conflict_T_9 = decode_entry_1_io_out_rs2 != 5'h0; // @[IDU.scala 184:34]
  wire  _self_reg_conflict_T_10 = (decode_entry_1_io_out_src2 == 2'h2 | decode_entry_1_io_out_fu_type == 3'h2) &
    _self_reg_conflict_T_9; // @[IDU.scala 183:92]
  wire  _self_reg_conflict_T_11 = decode_entry_1_io_out_rs2 == decode_entry_0_io_out_dest; // @[IDU.scala 185:34]
  wire  _self_reg_conflict_T_12 = _self_reg_conflict_T_10 & _self_reg_conflict_T_11; // @[IDU.scala 184:42]
  wire  _self_reg_conflict_T_13 = _self_reg_conflict_T_12 & decode_entry_0_io_out_wen; // @[IDU.scala 185:66]
  wire  self_reg_conflict = _self_reg_conflict_T_5 | _self_reg_conflict_T_13; // @[IDU.scala 182:33]
  wire  _self_fu_conflict_T_3 = decode_entry_0_io_out_fu_type == 3'h0 & decode_entry_1_io_out_fu_type == 3'h0; // @[IDU.scala 189:48]
  wire  self_fu_conflict = ~(decode_entry_0_io_out_fu_type != decode_entry_1_io_out_fu_type | _self_fu_conflict_T_3); // @[IDU.scala 188:23]
  wire  bpu_csr_conflict = decode_entry_0_io_out_fu_type == 3'h1 | decode_entry_0_io_out_fu_type == 3'h3 |
    decode_entry_1_io_out_fu_type == 3'h3; // @[IDU.scala 191:110]
  wire  _conflict_T_5 = self_fu_conflict | self_reg_conflict | bpu_csr_conflict; // @[IDU.scala 194:44]
  wire  conflict = decode_entry_1_io_out_valid & decode_entry_0_io_out_valid & io_in_valid & ~had_conflict &
    _conflict_T_5; // @[IDU.scala 193:110]
  wire  _io_out_bits_1_valid_T = ~conflict; // @[IDU.scala 196:59]
  wire  _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_20 = _T & conflict | had_conflict; // @[IDU.scala 198:34 IDU.scala 200:18 IDU.scala 174:29]
  wire  _GEN_41 = _T & had_conflict ? conflict_decode_entry_valid : decode_entry_0_io_out_valid; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  wire  _GEN_42 = _T & had_conflict ? 1'h0 : decode_entry_1_io_out_valid & ~conflict; // @[IDU.scala 203:38 IDU.scala 206:26 IDU.scala 196:24]
  Decode_Entry decode_entry_0 ( // @[IDU.scala 163:30]
    .io_in_valid(decode_entry_0_io_in_valid),
    .io_in_pc(decode_entry_0_io_in_pc),
    .io_in_inst(decode_entry_0_io_in_inst),
    .io_in_bp_br_taken(decode_entry_0_io_in_bp_br_taken),
    .io_in_bp_br_target(decode_entry_0_io_in_bp_br_target),
    .io_in_bp_br_type(decode_entry_0_io_in_bp_br_type),
    .io_out_valid(decode_entry_0_io_out_valid),
    .io_out_pc(decode_entry_0_io_out_pc),
    .io_out_inst(decode_entry_0_io_out_inst),
    .io_out_src1(decode_entry_0_io_out_src1),
    .io_out_src2(decode_entry_0_io_out_src2),
    .io_out_rs1(decode_entry_0_io_out_rs1),
    .io_out_rs2(decode_entry_0_io_out_rs2),
    .io_out_dest(decode_entry_0_io_out_dest),
    .io_out_imm(decode_entry_0_io_out_imm),
    .io_out_fu_type(decode_entry_0_io_out_fu_type),
    .io_out_bru_op(decode_entry_0_io_out_bru_op),
    .io_out_alu_op(decode_entry_0_io_out_alu_op),
    .io_out_lsu_op(decode_entry_0_io_out_lsu_op),
    .io_out_csr_op(decode_entry_0_io_out_csr_op),
    .io_out_mdu_op(decode_entry_0_io_out_mdu_op),
    .io_out_wen(decode_entry_0_io_out_wen),
    .io_out_rv64(decode_entry_0_io_out_rv64),
    .io_out_bp_br_taken(decode_entry_0_io_out_bp_br_taken),
    .io_out_bp_br_target(decode_entry_0_io_out_bp_br_target),
    .io_out_bp_br_type(decode_entry_0_io_out_bp_br_type)
  );
  Decode_Entry decode_entry_1 ( // @[IDU.scala 163:30]
    .io_in_valid(decode_entry_1_io_in_valid),
    .io_in_pc(decode_entry_1_io_in_pc),
    .io_in_inst(decode_entry_1_io_in_inst),
    .io_in_bp_br_taken(decode_entry_1_io_in_bp_br_taken),
    .io_in_bp_br_target(decode_entry_1_io_in_bp_br_target),
    .io_in_bp_br_type(decode_entry_1_io_in_bp_br_type),
    .io_out_valid(decode_entry_1_io_out_valid),
    .io_out_pc(decode_entry_1_io_out_pc),
    .io_out_inst(decode_entry_1_io_out_inst),
    .io_out_src1(decode_entry_1_io_out_src1),
    .io_out_src2(decode_entry_1_io_out_src2),
    .io_out_rs1(decode_entry_1_io_out_rs1),
    .io_out_rs2(decode_entry_1_io_out_rs2),
    .io_out_dest(decode_entry_1_io_out_dest),
    .io_out_imm(decode_entry_1_io_out_imm),
    .io_out_fu_type(decode_entry_1_io_out_fu_type),
    .io_out_bru_op(decode_entry_1_io_out_bru_op),
    .io_out_alu_op(decode_entry_1_io_out_alu_op),
    .io_out_lsu_op(decode_entry_1_io_out_lsu_op),
    .io_out_csr_op(decode_entry_1_io_out_csr_op),
    .io_out_mdu_op(decode_entry_1_io_out_mdu_op),
    .io_out_wen(decode_entry_1_io_out_wen),
    .io_out_rv64(decode_entry_1_io_out_rv64),
    .io_out_bp_br_taken(decode_entry_1_io_out_bp_br_taken),
    .io_out_bp_br_target(decode_entry_1_io_out_bp_br_target),
    .io_out_bp_br_type(decode_entry_1_io_out_bp_br_type)
  );
  assign io_in_ready = (io_out_ready | ~io_in_valid) & _io_out_bits_1_valid_T; // @[IDU.scala 219:49]
  assign io_out_valid = (io_in_valid | had_conflict) & ~frontend_reflush; // @[IDU.scala 218:49]
  assign io_out_bits_0_valid = frontend_reflush ? 1'h0 : _GEN_41; // @[IDU.scala 212:21 IDU.scala 214:26]
  assign io_out_bits_0_pc = _T & had_conflict ? conflict_decode_entry_pc : decode_entry_0_io_out_pc; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_inst = _T & had_conflict ? conflict_decode_entry_inst : decode_entry_0_io_out_inst; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_src1 = _T & had_conflict ? conflict_decode_entry_src1 : decode_entry_0_io_out_src1; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_src2 = _T & had_conflict ? conflict_decode_entry_src2 : decode_entry_0_io_out_src2; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_rs1 = _T & had_conflict ? conflict_decode_entry_rs1 : decode_entry_0_io_out_rs1; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_rs2 = _T & had_conflict ? conflict_decode_entry_rs2 : decode_entry_0_io_out_rs2; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_dest = _T & had_conflict ? conflict_decode_entry_dest : decode_entry_0_io_out_dest; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_imm = _T & had_conflict ? conflict_decode_entry_imm : decode_entry_0_io_out_imm; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_fu_type = _T & had_conflict ? conflict_decode_entry_fu_type : decode_entry_0_io_out_fu_type; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_bru_op = _T & had_conflict ? conflict_decode_entry_bru_op : decode_entry_0_io_out_bru_op; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_alu_op = _T & had_conflict ? conflict_decode_entry_alu_op : decode_entry_0_io_out_alu_op; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_lsu_op = _T & had_conflict ? conflict_decode_entry_lsu_op : decode_entry_0_io_out_lsu_op; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_csr_op = _T & had_conflict ? conflict_decode_entry_csr_op : decode_entry_0_io_out_csr_op; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_mdu_op = _T & had_conflict ? conflict_decode_entry_mdu_op : decode_entry_0_io_out_mdu_op; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_wen = _T & had_conflict ? conflict_decode_entry_wen : decode_entry_0_io_out_wen; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_rv64 = _T & had_conflict ? conflict_decode_entry_rv64 : decode_entry_0_io_out_rv64; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_bp_br_taken = _T & had_conflict ? conflict_decode_entry_bp_br_taken :
    decode_entry_0_io_out_bp_br_taken; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_bp_br_target = _T & had_conflict ? conflict_decode_entry_bp_br_target :
    decode_entry_0_io_out_bp_br_target; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_0_bp_br_type = _T & had_conflict ? conflict_decode_entry_bp_br_type :
    decode_entry_0_io_out_bp_br_type; // @[IDU.scala 203:38 IDU.scala 205:20 IDU.scala 169:28]
  assign io_out_bits_1_valid = frontend_reflush ? 1'h0 : _GEN_42; // @[IDU.scala 212:21 IDU.scala 215:26]
  assign io_out_bits_1_pc = decode_entry_1_io_out_pc; // @[IDU.scala 169:28]
  assign io_out_bits_1_inst = decode_entry_1_io_out_inst; // @[IDU.scala 169:28]
  assign io_out_bits_1_src1 = decode_entry_1_io_out_src1; // @[IDU.scala 169:28]
  assign io_out_bits_1_src2 = decode_entry_1_io_out_src2; // @[IDU.scala 169:28]
  assign io_out_bits_1_rs1 = decode_entry_1_io_out_rs1; // @[IDU.scala 169:28]
  assign io_out_bits_1_rs2 = decode_entry_1_io_out_rs2; // @[IDU.scala 169:28]
  assign io_out_bits_1_dest = decode_entry_1_io_out_dest; // @[IDU.scala 169:28]
  assign io_out_bits_1_imm = decode_entry_1_io_out_imm; // @[IDU.scala 169:28]
  assign io_out_bits_1_fu_type = decode_entry_1_io_out_fu_type; // @[IDU.scala 169:28]
  assign io_out_bits_1_bru_op = decode_entry_1_io_out_bru_op; // @[IDU.scala 169:28]
  assign io_out_bits_1_alu_op = decode_entry_1_io_out_alu_op; // @[IDU.scala 169:28]
  assign io_out_bits_1_lsu_op = decode_entry_1_io_out_lsu_op; // @[IDU.scala 169:28]
  assign io_out_bits_1_csr_op = decode_entry_1_io_out_csr_op; // @[IDU.scala 169:28]
  assign io_out_bits_1_mdu_op = decode_entry_1_io_out_mdu_op; // @[IDU.scala 169:28]
  assign io_out_bits_1_wen = decode_entry_1_io_out_wen; // @[IDU.scala 169:28]
  assign io_out_bits_1_rv64 = decode_entry_1_io_out_rv64; // @[IDU.scala 169:28]
  assign io_out_bits_1_bp_br_taken = decode_entry_1_io_out_bp_br_taken; // @[IDU.scala 169:28]
  assign io_out_bits_1_bp_br_target = decode_entry_1_io_out_bp_br_target; // @[IDU.scala 169:28]
  assign io_out_bits_1_bp_br_type = decode_entry_1_io_out_bp_br_type; // @[IDU.scala 169:28]
  assign decode_entry_0_io_in_valid = io_in_bits_0_valid; // @[IDU.scala 168:27]
  assign decode_entry_0_io_in_pc = io_in_bits_0_pc; // @[IDU.scala 168:27]
  assign decode_entry_0_io_in_inst = io_in_bits_0_inst; // @[IDU.scala 168:27]
  assign decode_entry_0_io_in_bp_br_taken = io_in_bits_0_bp_br_taken; // @[IDU.scala 168:27]
  assign decode_entry_0_io_in_bp_br_target = io_in_bits_0_bp_br_target; // @[IDU.scala 168:27]
  assign decode_entry_0_io_in_bp_br_type = io_in_bits_0_bp_br_type; // @[IDU.scala 168:27]
  assign decode_entry_1_io_in_valid = io_in_bits_1_valid; // @[IDU.scala 168:27]
  assign decode_entry_1_io_in_pc = io_in_bits_1_pc; // @[IDU.scala 168:27]
  assign decode_entry_1_io_in_inst = io_in_bits_1_inst; // @[IDU.scala 168:27]
  assign decode_entry_1_io_in_bp_br_taken = io_in_bits_1_bp_br_taken; // @[IDU.scala 168:27]
  assign decode_entry_1_io_in_bp_br_target = io_in_bits_1_bp_br_target; // @[IDU.scala 168:27]
  assign decode_entry_1_io_in_bp_br_type = io_in_bits_1_bp_br_type; // @[IDU.scala 168:27]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_valid <= 1'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_valid <= decode_entry_1_io_out_valid; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_pc <= 32'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_pc <= decode_entry_1_io_out_pc; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_inst <= 32'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_inst <= decode_entry_1_io_out_inst; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_src1 <= 2'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_src1 <= decode_entry_1_io_out_src1; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_src2 <= 2'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_src2 <= decode_entry_1_io_out_src2; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_rs1 <= 5'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_rs1 <= decode_entry_1_io_out_rs1; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_rs2 <= 5'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_rs2 <= decode_entry_1_io_out_rs2; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_dest <= 5'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_dest <= decode_entry_1_io_out_dest; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_imm <= 64'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_imm <= decode_entry_1_io_out_imm; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_fu_type <= 3'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_fu_type <= decode_entry_1_io_out_fu_type; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_bru_op <= 4'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_bru_op <= decode_entry_1_io_out_bru_op; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_alu_op <= 5'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_alu_op <= decode_entry_1_io_out_alu_op; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_lsu_op <= 4'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_lsu_op <= decode_entry_1_io_out_lsu_op; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_csr_op <= 3'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_csr_op <= decode_entry_1_io_out_csr_op; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_mdu_op <= 4'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_mdu_op <= decode_entry_1_io_out_mdu_op; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_wen <= 1'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_wen <= decode_entry_1_io_out_wen; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_rv64 <= 1'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_rv64 <= decode_entry_1_io_out_rv64; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_bp_br_taken <= 1'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_bp_br_taken <= decode_entry_1_io_out_bp_br_taken; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_bp_br_target <= 32'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_bp_br_target <= decode_entry_1_io_out_bp_br_target; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 172:38]
      conflict_decode_entry_bp_br_type <= 2'h0; // @[IDU.scala 172:38]
    end else if (_T & conflict) begin // @[IDU.scala 198:34]
      conflict_decode_entry_bp_br_type <= decode_entry_1_io_out_bp_br_type; // @[IDU.scala 199:27]
    end
    if (reset) begin // @[IDU.scala 174:29]
      had_conflict <= 1'h0; // @[IDU.scala 174:29]
    end else if (frontend_reflush) begin // @[IDU.scala 212:21]
      had_conflict <= 1'h0; // @[IDU.scala 213:18]
    end else if (_T & had_conflict) begin // @[IDU.scala 203:38]
      had_conflict <= 1'h0; // @[IDU.scala 204:18]
    end else begin
      had_conflict <= _GEN_20;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  conflict_decode_entry_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  conflict_decode_entry_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  conflict_decode_entry_inst = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  conflict_decode_entry_src1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  conflict_decode_entry_src2 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  conflict_decode_entry_rs1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  conflict_decode_entry_rs2 = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  conflict_decode_entry_dest = _RAND_7[4:0];
  _RAND_8 = {2{`RANDOM}};
  conflict_decode_entry_imm = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  conflict_decode_entry_fu_type = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  conflict_decode_entry_bru_op = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  conflict_decode_entry_alu_op = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  conflict_decode_entry_lsu_op = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  conflict_decode_entry_csr_op = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  conflict_decode_entry_mdu_op = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  conflict_decode_entry_wen = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  conflict_decode_entry_rv64 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  conflict_decode_entry_bp_br_taken = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  conflict_decode_entry_bp_br_target = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  conflict_decode_entry_bp_br_type = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  had_conflict = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Issue_Entry(
  input         io_in_valid,
  input  [31:0] io_in_pc,
  input  [31:0] io_in_inst,
  input  [1:0]  io_in_src1,
  input  [1:0]  io_in_src2,
  input  [4:0]  io_in_rs1,
  input  [4:0]  io_in_dest,
  input  [63:0] io_in_imm,
  input  [2:0]  io_in_fu_type,
  input  [3:0]  io_in_bru_op,
  input  [4:0]  io_in_alu_op,
  input  [3:0]  io_in_lsu_op,
  input  [2:0]  io_in_csr_op,
  input  [3:0]  io_in_mdu_op,
  input         io_in_wen,
  input         io_in_rv64,
  input         io_in_bp_br_taken,
  input  [31:0] io_in_bp_br_target,
  input  [1:0]  io_in_bp_br_type,
  output        io_out_valid,
  output [31:0] io_out_pc,
  output [31:0] io_out_inst,
  output [63:0] io_out_src1_value,
  output [63:0] io_out_src2_value,
  output [63:0] io_out_rs2_value,
  output [63:0] io_out_imm,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_dest,
  output [2:0]  io_out_fu_type,
  output [3:0]  io_out_bru_op,
  output [4:0]  io_out_alu_op,
  output [3:0]  io_out_lsu_op,
  output [2:0]  io_out_csr_op,
  output [3:0]  io_out_mdu_op,
  output        io_out_wen,
  output        io_out_rv64,
  output        io_out_bp_br_taken,
  output [31:0] io_out_bp_br_target,
  output [1:0]  io_out_bp_br_type,
  input  [63:0] io_rs1_value,
  input  [63:0] io_rs2_value
);
  wire [63:0] _src1_value_T = {59'h0,io_in_rs1}; // @[Cat.scala 30:58]
  wire [31:0] _src1_value_T_2 = 2'h1 == io_in_src1 ? io_in_pc : 32'h0; // @[Mux.scala 80:57]
  wire [63:0] _src1_value_T_4 = 2'h2 == io_in_src1 ? io_rs1_value : {{32'd0}, _src1_value_T_2}; // @[Mux.scala 80:57]
  wire [63:0] _src2_value_T_1 = 2'h2 == io_in_src2 ? io_rs2_value : 64'h0; // @[Mux.scala 80:57]
  assign io_out_valid = io_in_valid; // @[Issue.scala 42:13]
  assign io_out_pc = io_in_pc; // @[Issue.scala 43:10]
  assign io_out_inst = io_in_inst; // @[Issue.scala 44:12]
  assign io_out_src1_value = 2'h3 == io_in_src1 ? _src1_value_T : _src1_value_T_4; // @[Mux.scala 80:57]
  assign io_out_src2_value = 2'h3 == io_in_src2 ? io_in_imm : _src2_value_T_1; // @[Mux.scala 80:57]
  assign io_out_rs2_value = io_rs2_value; // @[Issue.scala 47:17]
  assign io_out_imm = io_in_imm; // @[Issue.scala 48:11]
  assign io_out_rs1 = io_in_rs1; // @[Issue.scala 49:11]
  assign io_out_dest = io_in_dest; // @[Issue.scala 50:12]
  assign io_out_fu_type = io_in_fu_type; // @[Issue.scala 51:15]
  assign io_out_bru_op = io_in_bru_op; // @[Issue.scala 53:14]
  assign io_out_alu_op = io_in_alu_op; // @[Issue.scala 52:14]
  assign io_out_lsu_op = io_in_lsu_op; // @[Issue.scala 54:14]
  assign io_out_csr_op = io_in_csr_op; // @[Issue.scala 55:14]
  assign io_out_mdu_op = io_in_mdu_op; // @[Issue.scala 56:14]
  assign io_out_wen = io_in_wen; // @[Issue.scala 57:11]
  assign io_out_rv64 = io_in_rv64; // @[Issue.scala 58:12]
  assign io_out_bp_br_taken = io_in_bp_br_taken; // @[Issue.scala 59:19]
  assign io_out_bp_br_target = io_in_bp_br_target; // @[Issue.scala 60:20]
  assign io_out_bp_br_type = io_in_bp_br_type; // @[Issue.scala 61:18]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [4:0]  io_rf_bus_0_raddr1,
  input  [4:0]  io_rf_bus_0_raddr2,
  output [63:0] io_rf_bus_0_rdata1,
  output [63:0] io_rf_bus_0_rdata2,
  input  [4:0]  io_rf_bus_0_waddr,
  input  [63:0] io_rf_bus_0_wdata,
  input         io_rf_bus_0_wen,
  input  [4:0]  io_rf_bus_1_raddr1,
  input  [4:0]  io_rf_bus_1_raddr2,
  output [63:0] io_rf_bus_1_rdata1,
  output [63:0] io_rf_bus_1_rdata2,
  input  [4:0]  io_rf_bus_1_waddr,
  input  [63:0] io_rf_bus_1_wdata,
  input         io_rf_bus_1_wen
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] rf_0; // @[RegFile.scala 11:19]
  reg [63:0] rf_1; // @[RegFile.scala 11:19]
  reg [63:0] rf_2; // @[RegFile.scala 11:19]
  reg [63:0] rf_3; // @[RegFile.scala 11:19]
  reg [63:0] rf_4; // @[RegFile.scala 11:19]
  reg [63:0] rf_5; // @[RegFile.scala 11:19]
  reg [63:0] rf_6; // @[RegFile.scala 11:19]
  reg [63:0] rf_7; // @[RegFile.scala 11:19]
  reg [63:0] rf_8; // @[RegFile.scala 11:19]
  reg [63:0] rf_9; // @[RegFile.scala 11:19]
  reg [63:0] rf_10; // @[RegFile.scala 11:19]
  reg [63:0] rf_11; // @[RegFile.scala 11:19]
  reg [63:0] rf_12; // @[RegFile.scala 11:19]
  reg [63:0] rf_13; // @[RegFile.scala 11:19]
  reg [63:0] rf_14; // @[RegFile.scala 11:19]
  reg [63:0] rf_15; // @[RegFile.scala 11:19]
  reg [63:0] rf_16; // @[RegFile.scala 11:19]
  reg [63:0] rf_17; // @[RegFile.scala 11:19]
  reg [63:0] rf_18; // @[RegFile.scala 11:19]
  reg [63:0] rf_19; // @[RegFile.scala 11:19]
  reg [63:0] rf_20; // @[RegFile.scala 11:19]
  reg [63:0] rf_21; // @[RegFile.scala 11:19]
  reg [63:0] rf_22; // @[RegFile.scala 11:19]
  reg [63:0] rf_23; // @[RegFile.scala 11:19]
  reg [63:0] rf_24; // @[RegFile.scala 11:19]
  reg [63:0] rf_25; // @[RegFile.scala 11:19]
  reg [63:0] rf_26; // @[RegFile.scala 11:19]
  reg [63:0] rf_27; // @[RegFile.scala 11:19]
  reg [63:0] rf_28; // @[RegFile.scala 11:19]
  reg [63:0] rf_29; // @[RegFile.scala 11:19]
  reg [63:0] rf_30; // @[RegFile.scala 11:19]
  reg [63:0] rf_31; // @[RegFile.scala 11:19]
  wire [63:0] _GEN_0 = 5'h0 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_0; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_1 = 5'h1 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_1; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_2 = 5'h2 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_2; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_3 = 5'h3 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_3; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_4 = 5'h4 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_4; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_5 = 5'h5 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_5; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_6 = 5'h6 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_6; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_7 = 5'h7 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_7; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_8 = 5'h8 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_8; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_9 = 5'h9 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_9; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_10 = 5'ha == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_10; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_11 = 5'hb == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_11; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_12 = 5'hc == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_12; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_13 = 5'hd == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_13; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_14 = 5'he == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_14; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_15 = 5'hf == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_15; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_16 = 5'h10 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_16; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_17 = 5'h11 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_17; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_18 = 5'h12 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_18; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_19 = 5'h13 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_19; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_20 = 5'h14 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_20; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_21 = 5'h15 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_21; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_22 = 5'h16 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_22; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_23 = 5'h17 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_23; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_24 = 5'h18 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_24; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_25 = 5'h19 == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_25; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_26 = 5'h1a == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_26; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_27 = 5'h1b == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_27; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_28 = 5'h1c == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_28; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_29 = 5'h1d == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_29; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_30 = 5'h1e == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_30; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_31 = 5'h1f == io_rf_bus_0_waddr ? io_rf_bus_0_wdata : rf_31; // @[RegFile.scala 15:27 RegFile.scala 15:27 RegFile.scala 11:19]
  wire [63:0] _GEN_32 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_0 : rf_0; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_33 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_1 : rf_1; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_34 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_2 : rf_2; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_35 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_3 : rf_3; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_36 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_4 : rf_4; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_37 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_5 : rf_5; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_38 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_6 : rf_6; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_39 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_7 : rf_7; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_40 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_8 : rf_8; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_41 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_9 : rf_9; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_42 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_10 : rf_10; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_43 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_11 : rf_11; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_44 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_12 : rf_12; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_45 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_13 : rf_13; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_46 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_14 : rf_14; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_47 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_15 : rf_15; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_48 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_16 : rf_16; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_49 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_17 : rf_17; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_50 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_18 : rf_18; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_51 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_19 : rf_19; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_52 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_20 : rf_20; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_53 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_21 : rf_21; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_54 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_22 : rf_22; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_55 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_23 : rf_23; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_56 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_24 : rf_24; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_57 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_25 : rf_25; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_58 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_26 : rf_26; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_59 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_27 : rf_27; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_60 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_28 : rf_28; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_61 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_29 : rf_29; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_62 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_30 : rf_30; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_63 = io_rf_bus_0_wen & io_rf_bus_0_waddr != 5'h0 ? _GEN_31 : rf_31; // @[RegFile.scala 14:55 RegFile.scala 11:19]
  wire [63:0] _GEN_65 = 5'h1 == io_rf_bus_0_raddr1 ? rf_1 : rf_0; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_66 = 5'h2 == io_rf_bus_0_raddr1 ? rf_2 : _GEN_65; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_67 = 5'h3 == io_rf_bus_0_raddr1 ? rf_3 : _GEN_66; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_68 = 5'h4 == io_rf_bus_0_raddr1 ? rf_4 : _GEN_67; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_69 = 5'h5 == io_rf_bus_0_raddr1 ? rf_5 : _GEN_68; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_70 = 5'h6 == io_rf_bus_0_raddr1 ? rf_6 : _GEN_69; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_71 = 5'h7 == io_rf_bus_0_raddr1 ? rf_7 : _GEN_70; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_72 = 5'h8 == io_rf_bus_0_raddr1 ? rf_8 : _GEN_71; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_73 = 5'h9 == io_rf_bus_0_raddr1 ? rf_9 : _GEN_72; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_74 = 5'ha == io_rf_bus_0_raddr1 ? rf_10 : _GEN_73; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_75 = 5'hb == io_rf_bus_0_raddr1 ? rf_11 : _GEN_74; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_76 = 5'hc == io_rf_bus_0_raddr1 ? rf_12 : _GEN_75; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_77 = 5'hd == io_rf_bus_0_raddr1 ? rf_13 : _GEN_76; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_78 = 5'he == io_rf_bus_0_raddr1 ? rf_14 : _GEN_77; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_79 = 5'hf == io_rf_bus_0_raddr1 ? rf_15 : _GEN_78; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_80 = 5'h10 == io_rf_bus_0_raddr1 ? rf_16 : _GEN_79; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_81 = 5'h11 == io_rf_bus_0_raddr1 ? rf_17 : _GEN_80; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_82 = 5'h12 == io_rf_bus_0_raddr1 ? rf_18 : _GEN_81; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_83 = 5'h13 == io_rf_bus_0_raddr1 ? rf_19 : _GEN_82; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_84 = 5'h14 == io_rf_bus_0_raddr1 ? rf_20 : _GEN_83; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_85 = 5'h15 == io_rf_bus_0_raddr1 ? rf_21 : _GEN_84; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_86 = 5'h16 == io_rf_bus_0_raddr1 ? rf_22 : _GEN_85; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_87 = 5'h17 == io_rf_bus_0_raddr1 ? rf_23 : _GEN_86; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_88 = 5'h18 == io_rf_bus_0_raddr1 ? rf_24 : _GEN_87; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_89 = 5'h19 == io_rf_bus_0_raddr1 ? rf_25 : _GEN_88; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_90 = 5'h1a == io_rf_bus_0_raddr1 ? rf_26 : _GEN_89; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_91 = 5'h1b == io_rf_bus_0_raddr1 ? rf_27 : _GEN_90; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_92 = 5'h1c == io_rf_bus_0_raddr1 ? rf_28 : _GEN_91; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_93 = 5'h1d == io_rf_bus_0_raddr1 ? rf_29 : _GEN_92; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_94 = 5'h1e == io_rf_bus_0_raddr1 ? rf_30 : _GEN_93; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_95 = 5'h1f == io_rf_bus_0_raddr1 ? rf_31 : _GEN_94; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_97 = 5'h1 == io_rf_bus_0_raddr2 ? rf_1 : rf_0; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_98 = 5'h2 == io_rf_bus_0_raddr2 ? rf_2 : _GEN_97; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_99 = 5'h3 == io_rf_bus_0_raddr2 ? rf_3 : _GEN_98; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_100 = 5'h4 == io_rf_bus_0_raddr2 ? rf_4 : _GEN_99; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_101 = 5'h5 == io_rf_bus_0_raddr2 ? rf_5 : _GEN_100; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_102 = 5'h6 == io_rf_bus_0_raddr2 ? rf_6 : _GEN_101; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_103 = 5'h7 == io_rf_bus_0_raddr2 ? rf_7 : _GEN_102; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_104 = 5'h8 == io_rf_bus_0_raddr2 ? rf_8 : _GEN_103; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_105 = 5'h9 == io_rf_bus_0_raddr2 ? rf_9 : _GEN_104; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_106 = 5'ha == io_rf_bus_0_raddr2 ? rf_10 : _GEN_105; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_107 = 5'hb == io_rf_bus_0_raddr2 ? rf_11 : _GEN_106; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_108 = 5'hc == io_rf_bus_0_raddr2 ? rf_12 : _GEN_107; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_109 = 5'hd == io_rf_bus_0_raddr2 ? rf_13 : _GEN_108; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_110 = 5'he == io_rf_bus_0_raddr2 ? rf_14 : _GEN_109; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_111 = 5'hf == io_rf_bus_0_raddr2 ? rf_15 : _GEN_110; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_112 = 5'h10 == io_rf_bus_0_raddr2 ? rf_16 : _GEN_111; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_113 = 5'h11 == io_rf_bus_0_raddr2 ? rf_17 : _GEN_112; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_114 = 5'h12 == io_rf_bus_0_raddr2 ? rf_18 : _GEN_113; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_115 = 5'h13 == io_rf_bus_0_raddr2 ? rf_19 : _GEN_114; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_116 = 5'h14 == io_rf_bus_0_raddr2 ? rf_20 : _GEN_115; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_117 = 5'h15 == io_rf_bus_0_raddr2 ? rf_21 : _GEN_116; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_118 = 5'h16 == io_rf_bus_0_raddr2 ? rf_22 : _GEN_117; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_119 = 5'h17 == io_rf_bus_0_raddr2 ? rf_23 : _GEN_118; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_120 = 5'h18 == io_rf_bus_0_raddr2 ? rf_24 : _GEN_119; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_121 = 5'h19 == io_rf_bus_0_raddr2 ? rf_25 : _GEN_120; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_122 = 5'h1a == io_rf_bus_0_raddr2 ? rf_26 : _GEN_121; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_123 = 5'h1b == io_rf_bus_0_raddr2 ? rf_27 : _GEN_122; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_124 = 5'h1c == io_rf_bus_0_raddr2 ? rf_28 : _GEN_123; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_125 = 5'h1d == io_rf_bus_0_raddr2 ? rf_29 : _GEN_124; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_126 = 5'h1e == io_rf_bus_0_raddr2 ? rf_30 : _GEN_125; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_127 = 5'h1f == io_rf_bus_0_raddr2 ? rf_31 : _GEN_126; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_193 = 5'h1 == io_rf_bus_1_raddr1 ? rf_1 : rf_0; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_194 = 5'h2 == io_rf_bus_1_raddr1 ? rf_2 : _GEN_193; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_195 = 5'h3 == io_rf_bus_1_raddr1 ? rf_3 : _GEN_194; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_196 = 5'h4 == io_rf_bus_1_raddr1 ? rf_4 : _GEN_195; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_197 = 5'h5 == io_rf_bus_1_raddr1 ? rf_5 : _GEN_196; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_198 = 5'h6 == io_rf_bus_1_raddr1 ? rf_6 : _GEN_197; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_199 = 5'h7 == io_rf_bus_1_raddr1 ? rf_7 : _GEN_198; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_200 = 5'h8 == io_rf_bus_1_raddr1 ? rf_8 : _GEN_199; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_201 = 5'h9 == io_rf_bus_1_raddr1 ? rf_9 : _GEN_200; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_202 = 5'ha == io_rf_bus_1_raddr1 ? rf_10 : _GEN_201; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_203 = 5'hb == io_rf_bus_1_raddr1 ? rf_11 : _GEN_202; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_204 = 5'hc == io_rf_bus_1_raddr1 ? rf_12 : _GEN_203; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_205 = 5'hd == io_rf_bus_1_raddr1 ? rf_13 : _GEN_204; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_206 = 5'he == io_rf_bus_1_raddr1 ? rf_14 : _GEN_205; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_207 = 5'hf == io_rf_bus_1_raddr1 ? rf_15 : _GEN_206; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_208 = 5'h10 == io_rf_bus_1_raddr1 ? rf_16 : _GEN_207; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_209 = 5'h11 == io_rf_bus_1_raddr1 ? rf_17 : _GEN_208; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_210 = 5'h12 == io_rf_bus_1_raddr1 ? rf_18 : _GEN_209; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_211 = 5'h13 == io_rf_bus_1_raddr1 ? rf_19 : _GEN_210; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_212 = 5'h14 == io_rf_bus_1_raddr1 ? rf_20 : _GEN_211; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_213 = 5'h15 == io_rf_bus_1_raddr1 ? rf_21 : _GEN_212; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_214 = 5'h16 == io_rf_bus_1_raddr1 ? rf_22 : _GEN_213; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_215 = 5'h17 == io_rf_bus_1_raddr1 ? rf_23 : _GEN_214; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_216 = 5'h18 == io_rf_bus_1_raddr1 ? rf_24 : _GEN_215; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_217 = 5'h19 == io_rf_bus_1_raddr1 ? rf_25 : _GEN_216; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_218 = 5'h1a == io_rf_bus_1_raddr1 ? rf_26 : _GEN_217; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_219 = 5'h1b == io_rf_bus_1_raddr1 ? rf_27 : _GEN_218; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_220 = 5'h1c == io_rf_bus_1_raddr1 ? rf_28 : _GEN_219; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_221 = 5'h1d == io_rf_bus_1_raddr1 ? rf_29 : _GEN_220; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_222 = 5'h1e == io_rf_bus_1_raddr1 ? rf_30 : _GEN_221; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_223 = 5'h1f == io_rf_bus_1_raddr1 ? rf_31 : _GEN_222; // @[RegFile.scala 17:28 RegFile.scala 17:28]
  wire [63:0] _GEN_225 = 5'h1 == io_rf_bus_1_raddr2 ? rf_1 : rf_0; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_226 = 5'h2 == io_rf_bus_1_raddr2 ? rf_2 : _GEN_225; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_227 = 5'h3 == io_rf_bus_1_raddr2 ? rf_3 : _GEN_226; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_228 = 5'h4 == io_rf_bus_1_raddr2 ? rf_4 : _GEN_227; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_229 = 5'h5 == io_rf_bus_1_raddr2 ? rf_5 : _GEN_228; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_230 = 5'h6 == io_rf_bus_1_raddr2 ? rf_6 : _GEN_229; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_231 = 5'h7 == io_rf_bus_1_raddr2 ? rf_7 : _GEN_230; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_232 = 5'h8 == io_rf_bus_1_raddr2 ? rf_8 : _GEN_231; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_233 = 5'h9 == io_rf_bus_1_raddr2 ? rf_9 : _GEN_232; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_234 = 5'ha == io_rf_bus_1_raddr2 ? rf_10 : _GEN_233; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_235 = 5'hb == io_rf_bus_1_raddr2 ? rf_11 : _GEN_234; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_236 = 5'hc == io_rf_bus_1_raddr2 ? rf_12 : _GEN_235; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_237 = 5'hd == io_rf_bus_1_raddr2 ? rf_13 : _GEN_236; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_238 = 5'he == io_rf_bus_1_raddr2 ? rf_14 : _GEN_237; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_239 = 5'hf == io_rf_bus_1_raddr2 ? rf_15 : _GEN_238; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_240 = 5'h10 == io_rf_bus_1_raddr2 ? rf_16 : _GEN_239; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_241 = 5'h11 == io_rf_bus_1_raddr2 ? rf_17 : _GEN_240; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_242 = 5'h12 == io_rf_bus_1_raddr2 ? rf_18 : _GEN_241; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_243 = 5'h13 == io_rf_bus_1_raddr2 ? rf_19 : _GEN_242; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_244 = 5'h14 == io_rf_bus_1_raddr2 ? rf_20 : _GEN_243; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_245 = 5'h15 == io_rf_bus_1_raddr2 ? rf_21 : _GEN_244; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_246 = 5'h16 == io_rf_bus_1_raddr2 ? rf_22 : _GEN_245; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_247 = 5'h17 == io_rf_bus_1_raddr2 ? rf_23 : _GEN_246; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_248 = 5'h18 == io_rf_bus_1_raddr2 ? rf_24 : _GEN_247; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_249 = 5'h19 == io_rf_bus_1_raddr2 ? rf_25 : _GEN_248; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_250 = 5'h1a == io_rf_bus_1_raddr2 ? rf_26 : _GEN_249; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_251 = 5'h1b == io_rf_bus_1_raddr2 ? rf_27 : _GEN_250; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_252 = 5'h1c == io_rf_bus_1_raddr2 ? rf_28 : _GEN_251; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_253 = 5'h1d == io_rf_bus_1_raddr2 ? rf_29 : _GEN_252; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_254 = 5'h1e == io_rf_bus_1_raddr2 ? rf_30 : _GEN_253; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  wire [63:0] _GEN_255 = 5'h1f == io_rf_bus_1_raddr2 ? rf_31 : _GEN_254; // @[RegFile.scala 18:28 RegFile.scala 18:28]
  assign io_rf_bus_0_rdata1 = io_rf_bus_0_raddr1 != 5'h0 ? _GEN_95 : 64'h0; // @[RegFile.scala 17:28]
  assign io_rf_bus_0_rdata2 = io_rf_bus_0_raddr2 != 5'h0 ? _GEN_127 : 64'h0; // @[RegFile.scala 18:28]
  assign io_rf_bus_1_rdata1 = io_rf_bus_1_raddr1 != 5'h0 ? _GEN_223 : 64'h0; // @[RegFile.scala 17:28]
  assign io_rf_bus_1_rdata2 = io_rf_bus_1_raddr2 != 5'h0 ? _GEN_255 : 64'h0; // @[RegFile.scala 18:28]
  always @(posedge clock) begin
    if (reset) begin // @[RegFile.scala 11:19]
      rf_0 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h0 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_0 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_0 <= _GEN_32;
      end
    end else begin
      rf_0 <= _GEN_32;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_1 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_1 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_1 <= _GEN_33;
      end
    end else begin
      rf_1 <= _GEN_33;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_2 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h2 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_2 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_2 <= _GEN_34;
      end
    end else begin
      rf_2 <= _GEN_34;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_3 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h3 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_3 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_3 <= _GEN_35;
      end
    end else begin
      rf_3 <= _GEN_35;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_4 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h4 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_4 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_4 <= _GEN_36;
      end
    end else begin
      rf_4 <= _GEN_36;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_5 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h5 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_5 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_5 <= _GEN_37;
      end
    end else begin
      rf_5 <= _GEN_37;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_6 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h6 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_6 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_6 <= _GEN_38;
      end
    end else begin
      rf_6 <= _GEN_38;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_7 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h7 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_7 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_7 <= _GEN_39;
      end
    end else begin
      rf_7 <= _GEN_39;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_8 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h8 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_8 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_8 <= _GEN_40;
      end
    end else begin
      rf_8 <= _GEN_40;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_9 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h9 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_9 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_9 <= _GEN_41;
      end
    end else begin
      rf_9 <= _GEN_41;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_10 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'ha == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_10 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_10 <= _GEN_42;
      end
    end else begin
      rf_10 <= _GEN_42;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_11 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'hb == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_11 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_11 <= _GEN_43;
      end
    end else begin
      rf_11 <= _GEN_43;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_12 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'hc == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_12 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_12 <= _GEN_44;
      end
    end else begin
      rf_12 <= _GEN_44;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_13 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'hd == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_13 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_13 <= _GEN_45;
      end
    end else begin
      rf_13 <= _GEN_45;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_14 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'he == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_14 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_14 <= _GEN_46;
      end
    end else begin
      rf_14 <= _GEN_46;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_15 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'hf == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_15 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_15 <= _GEN_47;
      end
    end else begin
      rf_15 <= _GEN_47;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_16 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h10 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_16 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_16 <= _GEN_48;
      end
    end else begin
      rf_16 <= _GEN_48;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_17 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h11 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_17 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_17 <= _GEN_49;
      end
    end else begin
      rf_17 <= _GEN_49;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_18 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h12 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_18 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_18 <= _GEN_50;
      end
    end else begin
      rf_18 <= _GEN_50;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_19 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h13 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_19 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_19 <= _GEN_51;
      end
    end else begin
      rf_19 <= _GEN_51;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_20 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h14 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_20 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_20 <= _GEN_52;
      end
    end else begin
      rf_20 <= _GEN_52;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_21 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h15 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_21 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_21 <= _GEN_53;
      end
    end else begin
      rf_21 <= _GEN_53;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_22 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h16 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_22 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_22 <= _GEN_54;
      end
    end else begin
      rf_22 <= _GEN_54;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_23 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h17 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_23 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_23 <= _GEN_55;
      end
    end else begin
      rf_23 <= _GEN_55;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_24 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h18 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_24 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_24 <= _GEN_56;
      end
    end else begin
      rf_24 <= _GEN_56;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_25 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h19 == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_25 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_25 <= _GEN_57;
      end
    end else begin
      rf_25 <= _GEN_57;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_26 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1a == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_26 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_26 <= _GEN_58;
      end
    end else begin
      rf_26 <= _GEN_58;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_27 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1b == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_27 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_27 <= _GEN_59;
      end
    end else begin
      rf_27 <= _GEN_59;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_28 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1c == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_28 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_28 <= _GEN_60;
      end
    end else begin
      rf_28 <= _GEN_60;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_29 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1d == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_29 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_29 <= _GEN_61;
      end
    end else begin
      rf_29 <= _GEN_61;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_30 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1e == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_30 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_30 <= _GEN_62;
      end
    end else begin
      rf_30 <= _GEN_62;
    end
    if (reset) begin // @[RegFile.scala 11:19]
      rf_31 <= 64'h0; // @[RegFile.scala 11:19]
    end else if (io_rf_bus_1_wen & io_rf_bus_1_waddr != 5'h0) begin // @[RegFile.scala 14:55]
      if (5'h1f == io_rf_bus_1_waddr) begin // @[RegFile.scala 15:27]
        rf_31 <= io_rf_bus_1_wdata; // @[RegFile.scala 15:27]
      end else begin
        rf_31 <= _GEN_63;
      end
    end else begin
      rf_31 <= _GEN_63;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rf_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  rf_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  rf_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  rf_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  rf_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  rf_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  rf_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  rf_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  rf_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  rf_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  rf_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  rf_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  rf_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  rf_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  rf_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  rf_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  rf_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  rf_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  rf_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  rf_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  rf_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  rf_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  rf_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  rf_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  rf_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  rf_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  rf_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  rf_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  rf_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  rf_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  rf_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  rf_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Issue(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_0_valid,
  input  [31:0] io_in_bits_0_pc,
  input  [31:0] io_in_bits_0_inst,
  input  [1:0]  io_in_bits_0_src1,
  input  [1:0]  io_in_bits_0_src2,
  input  [4:0]  io_in_bits_0_rs1,
  input  [4:0]  io_in_bits_0_rs2,
  input  [4:0]  io_in_bits_0_dest,
  input  [63:0] io_in_bits_0_imm,
  input  [2:0]  io_in_bits_0_fu_type,
  input  [3:0]  io_in_bits_0_bru_op,
  input  [4:0]  io_in_bits_0_alu_op,
  input  [3:0]  io_in_bits_0_lsu_op,
  input  [2:0]  io_in_bits_0_csr_op,
  input  [3:0]  io_in_bits_0_mdu_op,
  input         io_in_bits_0_wen,
  input         io_in_bits_0_rv64,
  input         io_in_bits_0_bp_br_taken,
  input  [31:0] io_in_bits_0_bp_br_target,
  input  [1:0]  io_in_bits_0_bp_br_type,
  input         io_in_bits_1_valid,
  input  [31:0] io_in_bits_1_pc,
  input  [31:0] io_in_bits_1_inst,
  input  [1:0]  io_in_bits_1_src1,
  input  [1:0]  io_in_bits_1_src2,
  input  [4:0]  io_in_bits_1_rs1,
  input  [4:0]  io_in_bits_1_rs2,
  input  [4:0]  io_in_bits_1_dest,
  input  [63:0] io_in_bits_1_imm,
  input  [2:0]  io_in_bits_1_fu_type,
  input  [3:0]  io_in_bits_1_bru_op,
  input  [4:0]  io_in_bits_1_alu_op,
  input  [3:0]  io_in_bits_1_lsu_op,
  input  [2:0]  io_in_bits_1_csr_op,
  input  [3:0]  io_in_bits_1_mdu_op,
  input         io_in_bits_1_wen,
  input         io_in_bits_1_rv64,
  input         io_in_bits_1_bp_br_taken,
  input  [31:0] io_in_bits_1_bp_br_target,
  input  [1:0]  io_in_bits_1_bp_br_type,
  input         io_out_ready,
  output        io_out_valid,
  output        io_out_bits_0_valid,
  output [31:0] io_out_bits_0_pc,
  output [31:0] io_out_bits_0_inst,
  output [63:0] io_out_bits_0_src1_value,
  output [63:0] io_out_bits_0_src2_value,
  output [63:0] io_out_bits_0_rs2_value,
  output [63:0] io_out_bits_0_imm,
  output [4:0]  io_out_bits_0_rs1,
  output [4:0]  io_out_bits_0_dest,
  output [2:0]  io_out_bits_0_fu_type,
  output [3:0]  io_out_bits_0_bru_op,
  output [4:0]  io_out_bits_0_alu_op,
  output [3:0]  io_out_bits_0_lsu_op,
  output [2:0]  io_out_bits_0_csr_op,
  output [3:0]  io_out_bits_0_mdu_op,
  output        io_out_bits_0_wen,
  output        io_out_bits_0_rv64,
  output        io_out_bits_0_bp_br_taken,
  output [31:0] io_out_bits_0_bp_br_target,
  output [1:0]  io_out_bits_0_bp_br_type,
  output        io_out_bits_1_valid,
  output [31:0] io_out_bits_1_pc,
  output [31:0] io_out_bits_1_inst,
  output [63:0] io_out_bits_1_src1_value,
  output [63:0] io_out_bits_1_src2_value,
  output [63:0] io_out_bits_1_rs2_value,
  output [63:0] io_out_bits_1_imm,
  output [4:0]  io_out_bits_1_rs1,
  output [4:0]  io_out_bits_1_dest,
  output [2:0]  io_out_bits_1_fu_type,
  output [3:0]  io_out_bits_1_bru_op,
  output [4:0]  io_out_bits_1_alu_op,
  output [3:0]  io_out_bits_1_lsu_op,
  output [2:0]  io_out_bits_1_csr_op,
  output [3:0]  io_out_bits_1_mdu_op,
  output        io_out_bits_1_wen,
  output        io_out_bits_1_rv64,
  output        io_out_bits_1_bp_br_taken,
  output [31:0] io_out_bits_1_bp_br_target,
  output [1:0]  io_out_bits_1_bp_br_type,
  input         io_wb_bus_0_rf_wen,
  input  [4:0]  io_wb_bus_0_rf_waddr,
  input  [63:0] io_wb_bus_0_rf_wdata,
  input         io_wb_bus_1_rf_wen,
  input  [4:0]  io_wb_bus_1_rf_waddr,
  input  [63:0] io_wb_bus_1_rf_wdata,
  input         io_ex_fwd_0_blk_valid,
  input         io_ex_fwd_0_fwd_valid,
  input  [4:0]  io_ex_fwd_0_rf_waddr,
  input  [63:0] io_ex_fwd_0_rf_wdata,
  input         io_ex_fwd_1_blk_valid,
  input         io_ex_fwd_1_fwd_valid,
  input  [4:0]  io_ex_fwd_1_rf_waddr,
  input  [63:0] io_ex_fwd_1_rf_wdata,
  input         frontend_reflush
);
  wire  issue_entry_0_io_in_valid; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_0_io_in_pc; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_0_io_in_inst; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_0_io_in_src1; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_0_io_in_src2; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_0_io_in_rs1; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_0_io_in_dest; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_in_imm; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_0_io_in_fu_type; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_0_io_in_bru_op; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_0_io_in_alu_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_0_io_in_lsu_op; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_0_io_in_csr_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_0_io_in_mdu_op; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_in_wen; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_in_rv64; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_in_bp_br_taken; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_0_io_in_bp_br_target; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_0_io_in_bp_br_type; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_out_valid; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_0_io_out_pc; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_0_io_out_inst; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_out_src1_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_out_src2_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_out_rs2_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_out_imm; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_0_io_out_rs1; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_0_io_out_dest; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_0_io_out_fu_type; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_0_io_out_bru_op; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_0_io_out_alu_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_0_io_out_lsu_op; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_0_io_out_csr_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_0_io_out_mdu_op; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_out_wen; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_out_rv64; // @[Issue.scala 83:29]
  wire  issue_entry_0_io_out_bp_br_taken; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_0_io_out_bp_br_target; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_0_io_out_bp_br_type; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_rs1_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_0_io_rs2_value; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_in_valid; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_1_io_in_pc; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_1_io_in_inst; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_1_io_in_src1; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_1_io_in_src2; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_1_io_in_rs1; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_1_io_in_dest; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_in_imm; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_1_io_in_fu_type; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_1_io_in_bru_op; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_1_io_in_alu_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_1_io_in_lsu_op; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_1_io_in_csr_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_1_io_in_mdu_op; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_in_wen; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_in_rv64; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_in_bp_br_taken; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_1_io_in_bp_br_target; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_1_io_in_bp_br_type; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_out_valid; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_1_io_out_pc; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_1_io_out_inst; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_out_src1_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_out_src2_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_out_rs2_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_out_imm; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_1_io_out_rs1; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_1_io_out_dest; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_1_io_out_fu_type; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_1_io_out_bru_op; // @[Issue.scala 83:29]
  wire [4:0] issue_entry_1_io_out_alu_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_1_io_out_lsu_op; // @[Issue.scala 83:29]
  wire [2:0] issue_entry_1_io_out_csr_op; // @[Issue.scala 83:29]
  wire [3:0] issue_entry_1_io_out_mdu_op; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_out_wen; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_out_rv64; // @[Issue.scala 83:29]
  wire  issue_entry_1_io_out_bp_br_taken; // @[Issue.scala 83:29]
  wire [31:0] issue_entry_1_io_out_bp_br_target; // @[Issue.scala 83:29]
  wire [1:0] issue_entry_1_io_out_bp_br_type; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_rs1_value; // @[Issue.scala 83:29]
  wire [63:0] issue_entry_1_io_rs2_value; // @[Issue.scala 83:29]
  wire  rf_clock; // @[Issue.scala 94:18]
  wire  rf_reset; // @[Issue.scala 94:18]
  wire [4:0] rf_io_rf_bus_0_raddr1; // @[Issue.scala 94:18]
  wire [4:0] rf_io_rf_bus_0_raddr2; // @[Issue.scala 94:18]
  wire [63:0] rf_io_rf_bus_0_rdata1; // @[Issue.scala 94:18]
  wire [63:0] rf_io_rf_bus_0_rdata2; // @[Issue.scala 94:18]
  wire [4:0] rf_io_rf_bus_0_waddr; // @[Issue.scala 94:18]
  wire [63:0] rf_io_rf_bus_0_wdata; // @[Issue.scala 94:18]
  wire  rf_io_rf_bus_0_wen; // @[Issue.scala 94:18]
  wire [4:0] rf_io_rf_bus_1_raddr1; // @[Issue.scala 94:18]
  wire [4:0] rf_io_rf_bus_1_raddr2; // @[Issue.scala 94:18]
  wire [63:0] rf_io_rf_bus_1_rdata1; // @[Issue.scala 94:18]
  wire [63:0] rf_io_rf_bus_1_rdata2; // @[Issue.scala 94:18]
  wire [4:0] rf_io_rf_bus_1_waddr; // @[Issue.scala 94:18]
  wire [63:0] rf_io_rf_bus_1_wdata; // @[Issue.scala 94:18]
  wire  rf_io_rf_bus_1_wen; // @[Issue.scala 94:18]
  wire  _rs1_value_0_T = io_ex_fwd_1_rf_waddr == io_in_bits_0_rs1; // @[Issue.scala 112:73]
  wire  _rs1_value_0_T_2 = io_ex_fwd_0_rf_waddr == io_in_bits_0_rs1; // @[Issue.scala 113:59]
  wire [63:0] _rs1_value_0_T_8 = io_wb_bus_0_rf_wen & io_wb_bus_0_rf_waddr == io_in_bits_0_rs1 ? io_wb_bus_0_rf_wdata :
    rf_io_rf_bus_0_rdata1; // @[Issue.scala 115:14]
  wire [63:0] _rs1_value_0_T_9 = io_wb_bus_1_rf_wen & io_wb_bus_1_rf_waddr == io_in_bits_0_rs1 ? io_wb_bus_1_rf_wdata :
    _rs1_value_0_T_8; // @[Issue.scala 114:12]
  wire [63:0] _rs1_value_0_T_10 = io_ex_fwd_0_fwd_valid & io_ex_fwd_0_rf_waddr == io_in_bits_0_rs1 ?
    io_ex_fwd_0_rf_wdata : _rs1_value_0_T_9; // @[Issue.scala 113:10]
  wire  _rs2_value_0_T = io_ex_fwd_1_rf_waddr == io_in_bits_0_rs2; // @[Issue.scala 117:73]
  wire  _rs2_value_0_T_2 = io_ex_fwd_0_rf_waddr == io_in_bits_0_rs2; // @[Issue.scala 118:59]
  wire [63:0] _rs2_value_0_T_8 = io_wb_bus_0_rf_wen & io_wb_bus_0_rf_waddr == io_in_bits_0_rs2 ? io_wb_bus_0_rf_wdata :
    rf_io_rf_bus_0_rdata2; // @[Issue.scala 120:14]
  wire [63:0] _rs2_value_0_T_9 = io_wb_bus_1_rf_wen & io_wb_bus_1_rf_waddr == io_in_bits_0_rs2 ? io_wb_bus_1_rf_wdata :
    _rs2_value_0_T_8; // @[Issue.scala 119:12]
  wire [63:0] _rs2_value_0_T_10 = io_ex_fwd_0_fwd_valid & io_ex_fwd_0_rf_waddr == io_in_bits_0_rs2 ?
    io_ex_fwd_0_rf_wdata : _rs2_value_0_T_9; // @[Issue.scala 118:10]
  wire  _need_blk_0_T_1 = io_in_bits_0_src1 == 2'h2; // @[Issue.scala 122:112]
  wire  _need_blk_0_T_4 = io_in_bits_0_src2 == 2'h2; // @[Issue.scala 123:71]
  wire  _need_blk_0_T_5 = _rs2_value_0_T_2 & io_in_bits_0_src2 == 2'h2; // @[Issue.scala 123:48]
  wire  _need_blk_0_T_7 = io_ex_fwd_0_blk_valid & (_rs1_value_0_T_2 & io_in_bits_0_src1 == 2'h2 | _need_blk_0_T_5); // @[Issue.scala 122:44]
  wire  _need_blk_0_T_13 = _rs2_value_0_T & _need_blk_0_T_4; // @[Issue.scala 125:50]
  wire  _need_blk_0_T_15 = io_ex_fwd_1_blk_valid & (_rs1_value_0_T & _need_blk_0_T_1 | _need_blk_0_T_13); // @[Issue.scala 124:31]
  wire  need_blk_0 = _need_blk_0_T_7 | _need_blk_0_T_15; // @[Issue.scala 123:85]
  wire  _rs1_value_1_T = io_ex_fwd_1_rf_waddr == io_in_bits_1_rs1; // @[Issue.scala 112:73]
  wire  _rs1_value_1_T_2 = io_ex_fwd_0_rf_waddr == io_in_bits_1_rs1; // @[Issue.scala 113:59]
  wire [63:0] _rs1_value_1_T_8 = io_wb_bus_0_rf_wen & io_wb_bus_0_rf_waddr == io_in_bits_1_rs1 ? io_wb_bus_0_rf_wdata :
    rf_io_rf_bus_1_rdata1; // @[Issue.scala 115:14]
  wire [63:0] _rs1_value_1_T_9 = io_wb_bus_1_rf_wen & io_wb_bus_1_rf_waddr == io_in_bits_1_rs1 ? io_wb_bus_1_rf_wdata :
    _rs1_value_1_T_8; // @[Issue.scala 114:12]
  wire [63:0] _rs1_value_1_T_10 = io_ex_fwd_0_fwd_valid & io_ex_fwd_0_rf_waddr == io_in_bits_1_rs1 ?
    io_ex_fwd_0_rf_wdata : _rs1_value_1_T_9; // @[Issue.scala 113:10]
  wire  _rs2_value_1_T = io_ex_fwd_1_rf_waddr == io_in_bits_1_rs2; // @[Issue.scala 117:73]
  wire  _rs2_value_1_T_2 = io_ex_fwd_0_rf_waddr == io_in_bits_1_rs2; // @[Issue.scala 118:59]
  wire [63:0] _rs2_value_1_T_8 = io_wb_bus_0_rf_wen & io_wb_bus_0_rf_waddr == io_in_bits_1_rs2 ? io_wb_bus_0_rf_wdata :
    rf_io_rf_bus_1_rdata2; // @[Issue.scala 120:14]
  wire [63:0] _rs2_value_1_T_9 = io_wb_bus_1_rf_wen & io_wb_bus_1_rf_waddr == io_in_bits_1_rs2 ? io_wb_bus_1_rf_wdata :
    _rs2_value_1_T_8; // @[Issue.scala 119:12]
  wire [63:0] _rs2_value_1_T_10 = io_ex_fwd_0_fwd_valid & io_ex_fwd_0_rf_waddr == io_in_bits_1_rs2 ?
    io_ex_fwd_0_rf_wdata : _rs2_value_1_T_9; // @[Issue.scala 118:10]
  wire  _need_blk_1_T_1 = io_in_bits_1_src1 == 2'h2; // @[Issue.scala 122:112]
  wire  _need_blk_1_T_4 = io_in_bits_1_src2 == 2'h2; // @[Issue.scala 123:71]
  wire  _need_blk_1_T_5 = _rs2_value_1_T_2 & io_in_bits_1_src2 == 2'h2; // @[Issue.scala 123:48]
  wire  _need_blk_1_T_7 = io_ex_fwd_0_blk_valid & (_rs1_value_1_T_2 & io_in_bits_1_src1 == 2'h2 | _need_blk_1_T_5); // @[Issue.scala 122:44]
  wire  _need_blk_1_T_13 = _rs2_value_1_T & _need_blk_1_T_4; // @[Issue.scala 125:50]
  wire  _need_blk_1_T_15 = io_ex_fwd_1_blk_valid & (_rs1_value_1_T & _need_blk_1_T_1 | _need_blk_1_T_13); // @[Issue.scala 124:31]
  wire  need_blk_1 = _need_blk_1_T_7 | _need_blk_1_T_15; // @[Issue.scala 123:85]
  wire [1:0] _io_out_valid_T = {need_blk_0,need_blk_1}; // @[Cat.scala 30:58]
  wire  _io_out_valid_T_2 = ~(|_io_out_valid_T); // @[Issue.scala 131:34]
  Issue_Entry issue_entry_0 ( // @[Issue.scala 83:29]
    .io_in_valid(issue_entry_0_io_in_valid),
    .io_in_pc(issue_entry_0_io_in_pc),
    .io_in_inst(issue_entry_0_io_in_inst),
    .io_in_src1(issue_entry_0_io_in_src1),
    .io_in_src2(issue_entry_0_io_in_src2),
    .io_in_rs1(issue_entry_0_io_in_rs1),
    .io_in_dest(issue_entry_0_io_in_dest),
    .io_in_imm(issue_entry_0_io_in_imm),
    .io_in_fu_type(issue_entry_0_io_in_fu_type),
    .io_in_bru_op(issue_entry_0_io_in_bru_op),
    .io_in_alu_op(issue_entry_0_io_in_alu_op),
    .io_in_lsu_op(issue_entry_0_io_in_lsu_op),
    .io_in_csr_op(issue_entry_0_io_in_csr_op),
    .io_in_mdu_op(issue_entry_0_io_in_mdu_op),
    .io_in_wen(issue_entry_0_io_in_wen),
    .io_in_rv64(issue_entry_0_io_in_rv64),
    .io_in_bp_br_taken(issue_entry_0_io_in_bp_br_taken),
    .io_in_bp_br_target(issue_entry_0_io_in_bp_br_target),
    .io_in_bp_br_type(issue_entry_0_io_in_bp_br_type),
    .io_out_valid(issue_entry_0_io_out_valid),
    .io_out_pc(issue_entry_0_io_out_pc),
    .io_out_inst(issue_entry_0_io_out_inst),
    .io_out_src1_value(issue_entry_0_io_out_src1_value),
    .io_out_src2_value(issue_entry_0_io_out_src2_value),
    .io_out_rs2_value(issue_entry_0_io_out_rs2_value),
    .io_out_imm(issue_entry_0_io_out_imm),
    .io_out_rs1(issue_entry_0_io_out_rs1),
    .io_out_dest(issue_entry_0_io_out_dest),
    .io_out_fu_type(issue_entry_0_io_out_fu_type),
    .io_out_bru_op(issue_entry_0_io_out_bru_op),
    .io_out_alu_op(issue_entry_0_io_out_alu_op),
    .io_out_lsu_op(issue_entry_0_io_out_lsu_op),
    .io_out_csr_op(issue_entry_0_io_out_csr_op),
    .io_out_mdu_op(issue_entry_0_io_out_mdu_op),
    .io_out_wen(issue_entry_0_io_out_wen),
    .io_out_rv64(issue_entry_0_io_out_rv64),
    .io_out_bp_br_taken(issue_entry_0_io_out_bp_br_taken),
    .io_out_bp_br_target(issue_entry_0_io_out_bp_br_target),
    .io_out_bp_br_type(issue_entry_0_io_out_bp_br_type),
    .io_rs1_value(issue_entry_0_io_rs1_value),
    .io_rs2_value(issue_entry_0_io_rs2_value)
  );
  Issue_Entry issue_entry_1 ( // @[Issue.scala 83:29]
    .io_in_valid(issue_entry_1_io_in_valid),
    .io_in_pc(issue_entry_1_io_in_pc),
    .io_in_inst(issue_entry_1_io_in_inst),
    .io_in_src1(issue_entry_1_io_in_src1),
    .io_in_src2(issue_entry_1_io_in_src2),
    .io_in_rs1(issue_entry_1_io_in_rs1),
    .io_in_dest(issue_entry_1_io_in_dest),
    .io_in_imm(issue_entry_1_io_in_imm),
    .io_in_fu_type(issue_entry_1_io_in_fu_type),
    .io_in_bru_op(issue_entry_1_io_in_bru_op),
    .io_in_alu_op(issue_entry_1_io_in_alu_op),
    .io_in_lsu_op(issue_entry_1_io_in_lsu_op),
    .io_in_csr_op(issue_entry_1_io_in_csr_op),
    .io_in_mdu_op(issue_entry_1_io_in_mdu_op),
    .io_in_wen(issue_entry_1_io_in_wen),
    .io_in_rv64(issue_entry_1_io_in_rv64),
    .io_in_bp_br_taken(issue_entry_1_io_in_bp_br_taken),
    .io_in_bp_br_target(issue_entry_1_io_in_bp_br_target),
    .io_in_bp_br_type(issue_entry_1_io_in_bp_br_type),
    .io_out_valid(issue_entry_1_io_out_valid),
    .io_out_pc(issue_entry_1_io_out_pc),
    .io_out_inst(issue_entry_1_io_out_inst),
    .io_out_src1_value(issue_entry_1_io_out_src1_value),
    .io_out_src2_value(issue_entry_1_io_out_src2_value),
    .io_out_rs2_value(issue_entry_1_io_out_rs2_value),
    .io_out_imm(issue_entry_1_io_out_imm),
    .io_out_rs1(issue_entry_1_io_out_rs1),
    .io_out_dest(issue_entry_1_io_out_dest),
    .io_out_fu_type(issue_entry_1_io_out_fu_type),
    .io_out_bru_op(issue_entry_1_io_out_bru_op),
    .io_out_alu_op(issue_entry_1_io_out_alu_op),
    .io_out_lsu_op(issue_entry_1_io_out_lsu_op),
    .io_out_csr_op(issue_entry_1_io_out_csr_op),
    .io_out_mdu_op(issue_entry_1_io_out_mdu_op),
    .io_out_wen(issue_entry_1_io_out_wen),
    .io_out_rv64(issue_entry_1_io_out_rv64),
    .io_out_bp_br_taken(issue_entry_1_io_out_bp_br_taken),
    .io_out_bp_br_target(issue_entry_1_io_out_bp_br_target),
    .io_out_bp_br_type(issue_entry_1_io_out_bp_br_type),
    .io_rs1_value(issue_entry_1_io_rs1_value),
    .io_rs2_value(issue_entry_1_io_rs2_value)
  );
  RegFile rf ( // @[Issue.scala 94:18]
    .clock(rf_clock),
    .reset(rf_reset),
    .io_rf_bus_0_raddr1(rf_io_rf_bus_0_raddr1),
    .io_rf_bus_0_raddr2(rf_io_rf_bus_0_raddr2),
    .io_rf_bus_0_rdata1(rf_io_rf_bus_0_rdata1),
    .io_rf_bus_0_rdata2(rf_io_rf_bus_0_rdata2),
    .io_rf_bus_0_waddr(rf_io_rf_bus_0_waddr),
    .io_rf_bus_0_wdata(rf_io_rf_bus_0_wdata),
    .io_rf_bus_0_wen(rf_io_rf_bus_0_wen),
    .io_rf_bus_1_raddr1(rf_io_rf_bus_1_raddr1),
    .io_rf_bus_1_raddr2(rf_io_rf_bus_1_raddr2),
    .io_rf_bus_1_rdata1(rf_io_rf_bus_1_rdata1),
    .io_rf_bus_1_rdata2(rf_io_rf_bus_1_rdata2),
    .io_rf_bus_1_waddr(rf_io_rf_bus_1_waddr),
    .io_rf_bus_1_wdata(rf_io_rf_bus_1_wdata),
    .io_rf_bus_1_wen(rf_io_rf_bus_1_wen)
  );
  assign io_in_ready = io_out_ready & _io_out_valid_T_2 | ~io_in_valid; // @[Issue.scala 132:55]
  assign io_out_valid = io_in_valid & ~(|_io_out_valid_T) & ~frontend_reflush; // @[Issue.scala 131:53]
  assign io_out_bits_0_valid = issue_entry_0_io_out_valid; // @[Issue.scala 89:27]
  assign io_out_bits_0_pc = issue_entry_0_io_out_pc; // @[Issue.scala 89:27]
  assign io_out_bits_0_inst = issue_entry_0_io_out_inst; // @[Issue.scala 89:27]
  assign io_out_bits_0_src1_value = issue_entry_0_io_out_src1_value; // @[Issue.scala 89:27]
  assign io_out_bits_0_src2_value = issue_entry_0_io_out_src2_value; // @[Issue.scala 89:27]
  assign io_out_bits_0_rs2_value = issue_entry_0_io_out_rs2_value; // @[Issue.scala 89:27]
  assign io_out_bits_0_imm = issue_entry_0_io_out_imm; // @[Issue.scala 89:27]
  assign io_out_bits_0_rs1 = issue_entry_0_io_out_rs1; // @[Issue.scala 89:27]
  assign io_out_bits_0_dest = issue_entry_0_io_out_dest; // @[Issue.scala 89:27]
  assign io_out_bits_0_fu_type = issue_entry_0_io_out_fu_type; // @[Issue.scala 89:27]
  assign io_out_bits_0_bru_op = issue_entry_0_io_out_bru_op; // @[Issue.scala 89:27]
  assign io_out_bits_0_alu_op = issue_entry_0_io_out_alu_op; // @[Issue.scala 89:27]
  assign io_out_bits_0_lsu_op = issue_entry_0_io_out_lsu_op; // @[Issue.scala 89:27]
  assign io_out_bits_0_csr_op = issue_entry_0_io_out_csr_op; // @[Issue.scala 89:27]
  assign io_out_bits_0_mdu_op = issue_entry_0_io_out_mdu_op; // @[Issue.scala 89:27]
  assign io_out_bits_0_wen = issue_entry_0_io_out_wen; // @[Issue.scala 89:27]
  assign io_out_bits_0_rv64 = issue_entry_0_io_out_rv64; // @[Issue.scala 89:27]
  assign io_out_bits_0_bp_br_taken = issue_entry_0_io_out_bp_br_taken; // @[Issue.scala 89:27]
  assign io_out_bits_0_bp_br_target = issue_entry_0_io_out_bp_br_target; // @[Issue.scala 89:27]
  assign io_out_bits_0_bp_br_type = issue_entry_0_io_out_bp_br_type; // @[Issue.scala 89:27]
  assign io_out_bits_1_valid = issue_entry_1_io_out_valid; // @[Issue.scala 89:27]
  assign io_out_bits_1_pc = issue_entry_1_io_out_pc; // @[Issue.scala 89:27]
  assign io_out_bits_1_inst = issue_entry_1_io_out_inst; // @[Issue.scala 89:27]
  assign io_out_bits_1_src1_value = issue_entry_1_io_out_src1_value; // @[Issue.scala 89:27]
  assign io_out_bits_1_src2_value = issue_entry_1_io_out_src2_value; // @[Issue.scala 89:27]
  assign io_out_bits_1_rs2_value = issue_entry_1_io_out_rs2_value; // @[Issue.scala 89:27]
  assign io_out_bits_1_imm = issue_entry_1_io_out_imm; // @[Issue.scala 89:27]
  assign io_out_bits_1_rs1 = issue_entry_1_io_out_rs1; // @[Issue.scala 89:27]
  assign io_out_bits_1_dest = issue_entry_1_io_out_dest; // @[Issue.scala 89:27]
  assign io_out_bits_1_fu_type = issue_entry_1_io_out_fu_type; // @[Issue.scala 89:27]
  assign io_out_bits_1_bru_op = issue_entry_1_io_out_bru_op; // @[Issue.scala 89:27]
  assign io_out_bits_1_alu_op = issue_entry_1_io_out_alu_op; // @[Issue.scala 89:27]
  assign io_out_bits_1_lsu_op = issue_entry_1_io_out_lsu_op; // @[Issue.scala 89:27]
  assign io_out_bits_1_csr_op = issue_entry_1_io_out_csr_op; // @[Issue.scala 89:27]
  assign io_out_bits_1_mdu_op = issue_entry_1_io_out_mdu_op; // @[Issue.scala 89:27]
  assign io_out_bits_1_wen = issue_entry_1_io_out_wen; // @[Issue.scala 89:27]
  assign io_out_bits_1_rv64 = issue_entry_1_io_out_rv64; // @[Issue.scala 89:27]
  assign io_out_bits_1_bp_br_taken = issue_entry_1_io_out_bp_br_taken; // @[Issue.scala 89:27]
  assign io_out_bits_1_bp_br_target = issue_entry_1_io_out_bp_br_target; // @[Issue.scala 89:27]
  assign io_out_bits_1_bp_br_type = issue_entry_1_io_out_bp_br_type; // @[Issue.scala 89:27]
  assign issue_entry_0_io_in_valid = io_in_bits_0_valid; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_pc = io_in_bits_0_pc; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_inst = io_in_bits_0_inst; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_src1 = io_in_bits_0_src1; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_src2 = io_in_bits_0_src2; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_rs1 = io_in_bits_0_rs1; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_dest = io_in_bits_0_dest; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_imm = io_in_bits_0_imm; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_fu_type = io_in_bits_0_fu_type; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_bru_op = io_in_bits_0_bru_op; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_alu_op = io_in_bits_0_alu_op; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_lsu_op = io_in_bits_0_lsu_op; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_csr_op = io_in_bits_0_csr_op; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_mdu_op = io_in_bits_0_mdu_op; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_wen = io_in_bits_0_wen; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_rv64 = io_in_bits_0_rv64; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_bp_br_taken = io_in_bits_0_bp_br_taken; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_bp_br_target = io_in_bits_0_bp_br_target; // @[Issue.scala 88:26]
  assign issue_entry_0_io_in_bp_br_type = io_in_bits_0_bp_br_type; // @[Issue.scala 88:26]
  assign issue_entry_0_io_rs1_value = io_ex_fwd_1_fwd_valid & io_ex_fwd_1_rf_waddr == io_in_bits_0_rs1 ?
    io_ex_fwd_1_rf_wdata : _rs1_value_0_T_10; // @[Issue.scala 112:24]
  assign issue_entry_0_io_rs2_value = io_ex_fwd_1_fwd_valid & io_ex_fwd_1_rf_waddr == io_in_bits_0_rs2 ?
    io_ex_fwd_1_rf_wdata : _rs2_value_0_T_10; // @[Issue.scala 117:24]
  assign issue_entry_1_io_in_valid = io_in_bits_1_valid; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_pc = io_in_bits_1_pc; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_inst = io_in_bits_1_inst; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_src1 = io_in_bits_1_src1; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_src2 = io_in_bits_1_src2; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_rs1 = io_in_bits_1_rs1; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_dest = io_in_bits_1_dest; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_imm = io_in_bits_1_imm; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_fu_type = io_in_bits_1_fu_type; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_bru_op = io_in_bits_1_bru_op; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_alu_op = io_in_bits_1_alu_op; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_lsu_op = io_in_bits_1_lsu_op; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_csr_op = io_in_bits_1_csr_op; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_mdu_op = io_in_bits_1_mdu_op; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_wen = io_in_bits_1_wen; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_rv64 = io_in_bits_1_rv64; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_bp_br_taken = io_in_bits_1_bp_br_taken; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_bp_br_target = io_in_bits_1_bp_br_target; // @[Issue.scala 88:26]
  assign issue_entry_1_io_in_bp_br_type = io_in_bits_1_bp_br_type; // @[Issue.scala 88:26]
  assign issue_entry_1_io_rs1_value = io_ex_fwd_1_fwd_valid & io_ex_fwd_1_rf_waddr == io_in_bits_1_rs1 ?
    io_ex_fwd_1_rf_wdata : _rs1_value_1_T_10; // @[Issue.scala 112:24]
  assign issue_entry_1_io_rs2_value = io_ex_fwd_1_fwd_valid & io_ex_fwd_1_rf_waddr == io_in_bits_1_rs2 ?
    io_ex_fwd_1_rf_wdata : _rs2_value_1_T_10; // @[Issue.scala 117:24]
  assign rf_clock = clock;
  assign rf_reset = reset;
  assign rf_io_rf_bus_0_raddr1 = io_in_bits_0_rs1; // @[Issue.scala 96:25]
  assign rf_io_rf_bus_0_raddr2 = io_in_bits_0_rs2; // @[Issue.scala 97:25]
  assign rf_io_rf_bus_0_waddr = io_wb_bus_0_rf_waddr; // @[Issue.scala 98:24]
  assign rf_io_rf_bus_0_wdata = io_wb_bus_0_rf_wdata; // @[Issue.scala 99:24]
  assign rf_io_rf_bus_0_wen = io_wb_bus_0_rf_wen; // @[Issue.scala 100:22]
  assign rf_io_rf_bus_1_raddr1 = io_in_bits_1_rs1; // @[Issue.scala 96:25]
  assign rf_io_rf_bus_1_raddr2 = io_in_bits_1_rs2; // @[Issue.scala 97:25]
  assign rf_io_rf_bus_1_waddr = io_wb_bus_1_rf_waddr; // @[Issue.scala 98:24]
  assign rf_io_rf_bus_1_wdata = io_wb_bus_1_rf_wdata; // @[Issue.scala 99:24]
  assign rf_io_rf_bus_1_wen = io_wb_bus_1_rf_wen; // @[Issue.scala 100:22]
endmodule
module ALU(
  input  [4:0]  io_alu_op,
  input         io_rv64,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  output [63:0] io_result
);
  wire  srl = io_alu_op == 5'h9 & io_rv64; // @[ALU.scala 19:31]
  wire  sra = io_alu_op == 5'ha & io_rv64; // @[ALU.scala 20:31]
  wire [31:0] src1_lo = io_src1[31:0]; // @[ALU.scala 23:38]
  wire [63:0] _src1_T = {32'h0,src1_lo}; // @[Cat.scala 30:58]
  wire [31:0] src1_hi_1 = io_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _src1_T_3 = {src1_hi_1,src1_lo}; // @[Cat.scala 30:58]
  wire [63:0] _src1_T_4 = sra ? _src1_T_3 : io_src1; // @[Mux.scala 98:16]
  wire [63:0] src1 = srl ? _src1_T : _src1_T_4; // @[Mux.scala 98:16]
  wire [5:0] shamt = io_rv64 ? {{1'd0}, io_src2[4:0]} : io_src2[5:0]; // @[ALU.scala 28:18]
  wire [63:0] _tmp_result_T_1 = src1 + io_src2; // @[ALU.scala 32:26]
  wire [63:0] _tmp_result_T_3 = src1 - io_src2; // @[ALU.scala 33:26]
  wire [63:0] _tmp_result_T_4 = src1 & io_src2; // @[ALU.scala 34:26]
  wire [63:0] _tmp_result_T_5 = src1 | io_src2; // @[ALU.scala 35:26]
  wire [63:0] _tmp_result_T_6 = src1 ^ io_src2; // @[ALU.scala 36:26]
  wire [63:0] _tmp_result_T_7 = srl ? _src1_T : _src1_T_4; // @[ALU.scala 37:26]
  wire  _tmp_result_T_9 = $signed(_tmp_result_T_7) < $signed(io_src2); // @[ALU.scala 37:33]
  wire  _tmp_result_T_10 = src1 < io_src2; // @[ALU.scala 38:26]
  wire [126:0] _GEN_0 = {{63'd0}, src1}; // @[ALU.scala 39:26]
  wire [126:0] _tmp_result_T_11 = _GEN_0 << shamt; // @[ALU.scala 39:26]
  wire [63:0] _tmp_result_T_12 = src1 >> shamt; // @[ALU.scala 40:26]
  wire [63:0] _tmp_result_T_15 = $signed(_tmp_result_T_7) >>> shamt; // @[ALU.scala 41:43]
  wire [63:0] _tmp_result_T_17 = 5'h1 == io_alu_op ? _tmp_result_T_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_19 = 5'h2 == io_alu_op ? _tmp_result_T_3 : _tmp_result_T_17; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_21 = 5'h3 == io_alu_op ? _tmp_result_T_4 : _tmp_result_T_19; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_23 = 5'h4 == io_alu_op ? _tmp_result_T_5 : _tmp_result_T_21; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_25 = 5'h5 == io_alu_op ? _tmp_result_T_6 : _tmp_result_T_23; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_27 = 5'h6 == io_alu_op ? {{63'd0}, _tmp_result_T_9} : _tmp_result_T_25; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_29 = 5'h7 == io_alu_op ? {{63'd0}, _tmp_result_T_10} : _tmp_result_T_27; // @[Mux.scala 80:57]
  wire [126:0] _tmp_result_T_31 = 5'h8 == io_alu_op ? _tmp_result_T_11 : {{63'd0}, _tmp_result_T_29}; // @[Mux.scala 80:57]
  wire [126:0] _tmp_result_T_33 = 5'h9 == io_alu_op ? {{63'd0}, _tmp_result_T_12} : _tmp_result_T_31; // @[Mux.scala 80:57]
  wire [126:0] _tmp_result_T_35 = 5'ha == io_alu_op ? {{63'd0}, _tmp_result_T_15} : _tmp_result_T_33; // @[Mux.scala 80:57]
  wire [63:0] tmp_result = _tmp_result_T_35[63:0]; // @[ALU.scala 29:24 ALU.scala 31:14]
  wire [31:0] io_result_hi = tmp_result[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_result_lo = tmp_result[31:0]; // @[ALU.scala 44:66]
  wire [63:0] _io_result_T_2 = {io_result_hi,io_result_lo}; // @[Cat.scala 30:58]
  assign io_result = io_rv64 ? _io_result_T_2 : tmp_result; // @[ALU.scala 44:19]
endmodule
module MDU(
  input         clock,
  input         reset,
  input  [3:0]  io_mdu_op,
  input         io_rv64,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  output        io_result_ok,
  output [63:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  src1_is_neg = io_src1[63]; // @[MDU.scala 20:25]
  wire  src2_is_neg = io_src2[63]; // @[MDU.scala 21:25]
  wire [63:0] _src1_abs_T = ~io_src1; // @[MDU.scala 22:36]
  wire [63:0] _src1_abs_T_2 = _src1_abs_T + 64'h1; // @[MDU.scala 22:50]
  wire [63:0] src1_abs = src1_is_neg ? _src1_abs_T_2 : io_src1; // @[MDU.scala 22:21]
  wire [63:0] _src2_abs_T = ~io_src2; // @[MDU.scala 23:36]
  wire [63:0] _src2_abs_T_2 = _src2_abs_T + 64'h1; // @[MDU.scala 23:50]
  wire [63:0] src2_abs = src2_is_neg ? _src2_abs_T_2 : io_src2; // @[MDU.scala 23:21]
  wire  is_mul = io_mdu_op == 4'h1 | io_mdu_op == 4'h2 | io_mdu_op == 4'h3 | io_mdu_op == 4'h4; // @[MDU.scala 27:89]
  wire  is_div = io_mdu_op == 4'h5 | io_mdu_op == 4'h6 | io_mdu_op == 4'h7 | io_mdu_op == 4'h8; // @[MDU.scala 28:86]
  wire  _src1_need_neg_T_5 = 4'h3 == io_mdu_op ? src1_is_neg : 4'h2 == io_mdu_op & src1_is_neg; // @[Mux.scala 80:57]
  wire  _src1_need_neg_T_7 = 4'h4 == io_mdu_op ? 1'h0 : _src1_need_neg_T_5; // @[Mux.scala 80:57]
  wire  _src1_need_neg_T_9 = 4'h5 == io_mdu_op ? src1_is_neg : _src1_need_neg_T_7; // @[Mux.scala 80:57]
  wire  _src1_need_neg_T_11 = 4'h6 == io_mdu_op ? 1'h0 : _src1_need_neg_T_9; // @[Mux.scala 80:57]
  wire  _src1_need_neg_T_13 = 4'h7 == io_mdu_op ? src1_is_neg : _src1_need_neg_T_11; // @[Mux.scala 80:57]
  wire  src1_need_neg = 4'h8 == io_mdu_op ? 1'h0 : _src1_need_neg_T_13; // @[Mux.scala 80:57]
  wire [63:0] src1_final = src1_need_neg ? src1_abs : io_src1; // @[MDU.scala 29:23]
  wire [63:0] src2_final = src1_need_neg ? src2_abs : io_src2; // @[MDU.scala 30:23]
  wire  _src2_need_neg_T_5 = 4'h3 == io_mdu_op ? 1'h0 : 4'h2 == io_mdu_op & src2_is_neg; // @[Mux.scala 80:57]
  wire  _src2_need_neg_T_7 = 4'h4 == io_mdu_op ? 1'h0 : _src2_need_neg_T_5; // @[Mux.scala 80:57]
  wire  _src2_need_neg_T_9 = 4'h5 == io_mdu_op ? src2_is_neg : _src2_need_neg_T_7; // @[Mux.scala 80:57]
  wire  _src2_need_neg_T_11 = 4'h6 == io_mdu_op ? 1'h0 : _src2_need_neg_T_9; // @[Mux.scala 80:57]
  wire  _src2_need_neg_T_13 = 4'h7 == io_mdu_op ? src2_is_neg : _src2_need_neg_T_11; // @[Mux.scala 80:57]
  wire  src2_need_neg = 4'h8 == io_mdu_op ? 1'h0 : _src2_need_neg_T_13; // @[Mux.scala 80:57]
  wire  result_is_neg = src1_need_neg ^ src2_need_neg; // @[LFSR.scala 15:41]
  reg [1:0] state; // @[MDU.scala 58:22]
  reg [5:0] count; // @[MDU.scala 59:22]
  wire [5:0] count_reverse = 6'h3f - count; // @[MDU.scala 60:28]
  reg [127:0] result_reg; // @[MDU.scala 61:27]
  reg [127:0] divisor_reg; // @[MDU.scala 62:28]
  reg [63:0] div_result_reg; // @[MDU.scala 63:31]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [127:0] _result_reg_T = {64'h0,src1_final}; // @[Cat.scala 30:58]
  wire [128:0] _result_reg_T_1 = {_result_reg_T, 1'h0}; // @[MDU.scala 73:54]
  wire [127:0] _divisor_reg_T = {src2_final,64'h0}; // @[Cat.scala 30:58]
  wire [128:0] _GEN_1 = is_div ? _result_reg_T_1 : {{1'd0}, result_reg}; // @[MDU.scala 71:28 MDU.scala 73:20 MDU.scala 61:27]
  wire [63:0] _GEN_3 = is_div ? 64'h0 : div_result_reg; // @[MDU.scala 71:28 MDU.scala 75:24 MDU.scala 63:31]
  wire [128:0] _GEN_5 = is_mul ? 129'h0 : _GEN_1; // @[MDU.scala 68:21 MDU.scala 70:20]
  wire [63:0] _GEN_7 = is_mul ? div_result_reg : _GEN_3; // @[MDU.scala 68:21 MDU.scala 63:31]
  wire  _T_1 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [63:0] _T_2 = src2_final >> count_reverse; // @[MDU.scala 79:23]
  wire [128:0] _result_reg_T_2 = {result_reg, 1'h0}; // @[MDU.scala 80:35]
  wire [128:0] _GEN_34 = {{65'd0}, src1_final}; // @[MDU.scala 80:50]
  wire [128:0] _result_reg_T_4 = _result_reg_T_2 + _GEN_34; // @[MDU.scala 80:50]
  wire [128:0] _GEN_8 = _T_2[0] ? _result_reg_T_4 : _result_reg_T_2; // @[MDU.scala 79:48 MDU.scala 80:20 MDU.scala 82:20]
  wire  _T_5 = count == 6'h3f; // @[MDU.scala 84:19]
  wire [5:0] _count_T_1 = count + 6'h1; // @[MDU.scala 87:24]
  wire [1:0] _GEN_9 = count == 6'h3f ? 2'h3 : state; // @[MDU.scala 84:29 MDU.scala 85:15 MDU.scala 58:22]
  wire [5:0] _GEN_10 = count == 6'h3f ? count : _count_T_1; // @[MDU.scala 84:29 MDU.scala 59:22 MDU.scala 87:15]
  wire  _T_6 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = result_reg[127:64] >= divisor_reg[127:64]; // @[MDU.scala 93:34]
  wire [127:0] _result_reg_T_7 = result_reg - divisor_reg; // @[MDU.scala 94:36]
  wire [64:0] _div_result_reg_T = {div_result_reg, 1'h0}; // @[MDU.scala 95:45]
  wire [64:0] _div_result_reg_T_2 = _div_result_reg_T + 65'h1; // @[MDU.scala 95:60]
  wire [127:0] _GEN_11 = result_reg[127:64] >= divisor_reg[127:64] ? _result_reg_T_7 : result_reg; // @[MDU.scala 93:59 MDU.scala 94:22 MDU.scala 61:27]
  wire [64:0] _GEN_12 = result_reg[127:64] >= divisor_reg[127:64] ? _div_result_reg_T_2 : _div_result_reg_T; // @[MDU.scala 93:59 MDU.scala 95:26 MDU.scala 97:26]
  wire [128:0] _result_reg_T_10 = {_result_reg_T_7, 1'h0}; // @[MDU.scala 102:52]
  wire [128:0] _GEN_13 = _T_10 ? _result_reg_T_10 : _result_reg_T_2; // @[MDU.scala 101:59 MDU.scala 102:22 MDU.scala 105:22]
  wire [128:0] _GEN_16 = _T_5 ? {{1'd0}, _GEN_11} : _GEN_13; // @[MDU.scala 91:29]
  wire [64:0] _GEN_17 = _T_5 ? _GEN_12 : _GEN_12; // @[MDU.scala 91:29]
  wire  _T_14 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_19 = _T_14 ? 2'h0 : state; // @[Conditional.scala 39:67 MDU.scala 111:13 MDU.scala 58:22]
  wire [5:0] _GEN_20 = _T_14 ? 6'h0 : count; // @[Conditional.scala 39:67 MDU.scala 112:13 MDU.scala 59:22]
  wire [128:0] _GEN_22 = _T_6 ? _GEN_16 : {{1'd0}, result_reg}; // @[Conditional.scala 39:67 MDU.scala 61:27]
  wire [64:0] _GEN_23 = _T_6 ? _GEN_17 : {{1'd0}, div_result_reg}; // @[Conditional.scala 39:67 MDU.scala 63:31]
  wire [128:0] _GEN_25 = _T_1 ? _GEN_8 : _GEN_22; // @[Conditional.scala 39:67]
  wire [64:0] _GEN_28 = _T_1 ? {{1'd0}, div_result_reg} : _GEN_23; // @[Conditional.scala 39:67 MDU.scala 63:31]
  wire [128:0] _GEN_30 = _T ? _GEN_5 : _GEN_25; // @[Conditional.scala 40:58]
  wire [64:0] _GEN_32 = _T ? {{1'd0}, _GEN_7} : _GEN_28; // @[Conditional.scala 40:58]
  wire [63:0] _tmp_result_T_1 = ~result_reg[63:0]; // @[MDU.scala 118:36]
  wire [63:0] _tmp_result_T_3 = _tmp_result_T_1 + 64'h1; // @[MDU.scala 118:63]
  wire [63:0] _tmp_result_T_5 = result_is_neg ? _tmp_result_T_3 : result_reg[63:0]; // @[MDU.scala 118:19]
  wire [63:0] _tmp_result_T_7 = ~result_reg[127:64]; // @[MDU.scala 119:37]
  wire [63:0] _tmp_result_T_9 = _tmp_result_T_7 + 64'h1; // @[MDU.scala 119:66]
  wire [63:0] _tmp_result_T_11 = result_is_neg ? _tmp_result_T_9 : result_reg[127:64]; // @[MDU.scala 119:20]
  wire [63:0] _tmp_result_T_24 = ~div_result_reg; // @[MDU.scala 122:36]
  wire [63:0] _tmp_result_T_26 = _tmp_result_T_24 + 64'h1; // @[MDU.scala 122:60]
  wire [63:0] _tmp_result_T_27 = result_is_neg ? _tmp_result_T_26 : div_result_reg; // @[MDU.scala 122:19]
  wire [63:0] _tmp_result_T_45 = 4'h1 == io_mdu_op ? _tmp_result_T_5 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_47 = 4'h2 == io_mdu_op ? _tmp_result_T_11 : _tmp_result_T_45; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_49 = 4'h3 == io_mdu_op ? _tmp_result_T_11 : _tmp_result_T_47; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_51 = 4'h4 == io_mdu_op ? _tmp_result_T_11 : _tmp_result_T_49; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_53 = 4'h5 == io_mdu_op ? _tmp_result_T_27 : _tmp_result_T_51; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_55 = 4'h6 == io_mdu_op ? _tmp_result_T_27 : _tmp_result_T_53; // @[Mux.scala 80:57]
  wire [63:0] _tmp_result_T_57 = 4'h7 == io_mdu_op ? _tmp_result_T_11 : _tmp_result_T_55; // @[Mux.scala 80:57]
  wire [63:0] tmp_result = 4'h8 == io_mdu_op ? _tmp_result_T_11 : _tmp_result_T_57; // @[Mux.scala 80:57]
  wire [31:0] io_result_hi = tmp_result[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] io_result_lo = tmp_result[31:0]; // @[MDU.scala 127:69]
  wire [63:0] _io_result_T_2 = {io_result_hi,io_result_lo}; // @[Cat.scala 30:58]
  assign io_result_ok = state == 2'h3; // @[MDU.scala 116:25]
  assign io_result = io_rv64 ? _io_result_T_2 : tmp_result; // @[MDU.scala 127:19]
  always @(posedge clock) begin
    if (reset) begin // @[MDU.scala 58:22]
      state <= 2'h0; // @[MDU.scala 58:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (is_mul) begin // @[MDU.scala 68:21]
        state <= 2'h1; // @[MDU.scala 69:15]
      end else if (is_div) begin // @[MDU.scala 71:28]
        state <= 2'h2; // @[MDU.scala 72:15]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      state <= _GEN_9;
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_9;
    end else begin
      state <= _GEN_19;
    end
    if (reset) begin // @[MDU.scala 59:22]
      count <= 6'h0; // @[MDU.scala 59:22]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        count <= _GEN_10;
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        count <= _GEN_10;
      end else begin
        count <= _GEN_20;
      end
    end
    if (reset) begin // @[MDU.scala 61:27]
      result_reg <= 128'h0; // @[MDU.scala 61:27]
    end else begin
      result_reg <= _GEN_30[127:0];
    end
    if (reset) begin // @[MDU.scala 62:28]
      divisor_reg <= 128'h0; // @[MDU.scala 62:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (!(is_mul)) begin // @[MDU.scala 68:21]
        if (is_div) begin // @[MDU.scala 71:28]
          divisor_reg <= _divisor_reg_T; // @[MDU.scala 74:21]
        end
      end
    end
    if (reset) begin // @[MDU.scala 63:31]
      div_result_reg <= 64'h0; // @[MDU.scala 63:31]
    end else begin
      div_result_reg <= _GEN_32[63:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  count = _RAND_1[5:0];
  _RAND_2 = {4{`RANDOM}};
  result_reg = _RAND_2[127:0];
  _RAND_3 = {4{`RANDOM}};
  divisor_reg = _RAND_3[127:0];
  _RAND_4 = {2{`RANDOM}};
  div_result_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BRU(
  input  [3:0]  io_bru_op,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [31:0] io_pc,
  input  [63:0] io_imm,
  output        io_br_taken,
  output [31:0] io_br_target,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rd,
  output [1:0]  io_btb_type
);
  wire  _io_br_taken_T = io_src1 == io_src2; // @[BRU.scala 26:26]
  wire  _io_br_taken_T_1 = io_src1 != io_src2; // @[BRU.scala 27:26]
  wire  _io_br_taken_T_4 = $signed(io_src1) < $signed(io_src2); // @[BRU.scala 28:33]
  wire  _io_br_taken_T_7 = $signed(io_src1) >= $signed(io_src2); // @[BRU.scala 29:33]
  wire  _io_br_taken_T_8 = io_src1 < io_src2; // @[BRU.scala 30:33]
  wire  _io_br_taken_T_9 = io_src1 >= io_src2; // @[BRU.scala 31:33]
  wire  _io_br_taken_T_15 = 4'h3 == io_bru_op ? _io_br_taken_T : 4'h2 == io_bru_op | 4'h1 == io_bru_op; // @[Mux.scala 80:57]
  wire  _io_br_taken_T_17 = 4'h4 == io_bru_op ? _io_br_taken_T_1 : _io_br_taken_T_15; // @[Mux.scala 80:57]
  wire  _io_br_taken_T_19 = 4'h5 == io_bru_op ? _io_br_taken_T_4 : _io_br_taken_T_17; // @[Mux.scala 80:57]
  wire  _io_br_taken_T_21 = 4'h6 == io_bru_op ? _io_br_taken_T_7 : _io_br_taken_T_19; // @[Mux.scala 80:57]
  wire  _io_br_taken_T_23 = 4'h7 == io_bru_op ? _io_br_taken_T_8 : _io_br_taken_T_21; // @[Mux.scala 80:57]
  wire  _io_br_target_T = io_bru_op == 4'h2; // @[BRU.scala 34:33]
  wire [31:0] _io_br_target_T_4 = io_src1[31:0] + io_imm[31:0]; // @[BRU.scala 34:64]
  wire [31:0] _io_br_target_T_6 = {_io_br_target_T_4[31:1], 1'h0}; // @[BRU.scala 34:87]
  wire [31:0] _io_br_target_T_10 = io_pc + io_imm[31:0]; // @[BRU.scala 34:106]
  wire  _T_2 = io_bru_op == 4'h1 | _io_br_target_T; // @[BRU.scala 36:32]
  wire [1:0] _GEN_0 = _T_2 ? 2'h3 : 2'h2; // @[BRU.scala 40:65 BRU.scala 41:14 BRU.scala 43:14]
  wire [1:0] _GEN_1 = _io_br_target_T & io_rs1 == 5'h1 ? 2'h1 : _GEN_0; // @[BRU.scala 38:60 BRU.scala 39:14]
  assign io_br_taken = 4'h8 == io_bru_op ? _io_br_taken_T_9 : _io_br_taken_T_23; // @[Mux.scala 80:57]
  assign io_br_target = io_bru_op == 4'h2 ? _io_br_target_T_6 : _io_br_target_T_10; // @[BRU.scala 34:22]
  assign io_btb_type = (io_bru_op == 4'h1 | _io_br_target_T) & io_rd == 5'h1 ? 2'h0 : _GEN_1; // @[BRU.scala 36:77 BRU.scala 37:14]
endmodule
module LSU(
  input         clock,
  input         reset,
  output        io_dmem_valid,
  output        io_dmem_op,
  output [31:0] io_dmem_addr,
  output [7:0]  io_dmem_wstrb,
  output [63:0] io_dmem_wdata,
  output        io_dmem_fence,
  input         io_dmem_fence_finish,
  input         io_dmem_data_ok,
  input  [63:0] io_dmem_rdata,
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [63:0] io_wdata,
  output [31:0] io_addr,
  input         io_is_lsu,
  input         io_wen,
  input  [3:0]  io_lsu_op,
  output [63:0] io_rdata,
  input         io_is_mdu,
  input         io_mdu_ok,
  output        dcache_fence_finish_0,
  input         fence_i,
  input         icache_fence_finish_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] _io_addr_T_1 = io_src1 + io_src2; // @[LSU.scala 28:23]
  wire [2:0] addr_low = io_addr[2:0]; // @[LSU.scala 29:22]
  wire [7:0] sb_wdata_hi = io_wdata[7:0]; // @[LSU.scala 53:28]
  wire [63:0] sb_wdata = {sb_wdata_hi,sb_wdata_hi,sb_wdata_hi,sb_wdata_hi,sb_wdata_hi,sb_wdata_hi,sb_wdata_hi,
    sb_wdata_hi}; // @[Cat.scala 30:58]
  wire [15:0] sh_wdata_hi = io_wdata[15:0]; // @[LSU.scala 54:28]
  wire [63:0] sh_wdata = {sh_wdata_hi,sh_wdata_hi,sh_wdata_hi,sh_wdata_hi}; // @[Cat.scala 30:58]
  wire [31:0] sw_wdata_hi = io_wdata[31:0]; // @[LSU.scala 55:28]
  wire [63:0] sw_wdata = {sw_wdata_hi,sw_wdata_hi}; // @[Cat.scala 30:58]
  wire [63:0] _dmem_wdata_T_1 = 4'h6 == io_lsu_op ? sb_wdata : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _dmem_wdata_T_3 = 4'h7 == io_lsu_op ? sh_wdata : _dmem_wdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _dmem_wdata_T_5 = 4'h8 == io_lsu_op ? sw_wdata : _dmem_wdata_T_3; // @[Mux.scala 80:57]
  wire [1:0] _sb_wmask_T_1 = 3'h1 == addr_low ? 2'h2 : 2'h1; // @[Mux.scala 80:57]
  wire [2:0] _sb_wmask_T_3 = 3'h2 == addr_low ? 3'h4 : {{1'd0}, _sb_wmask_T_1}; // @[Mux.scala 80:57]
  wire [3:0] _sb_wmask_T_5 = 3'h3 == addr_low ? 4'h8 : {{1'd0}, _sb_wmask_T_3}; // @[Mux.scala 80:57]
  wire [4:0] _sb_wmask_T_7 = 3'h4 == addr_low ? 5'h10 : {{1'd0}, _sb_wmask_T_5}; // @[Mux.scala 80:57]
  wire [5:0] _sb_wmask_T_9 = 3'h5 == addr_low ? 6'h20 : {{1'd0}, _sb_wmask_T_7}; // @[Mux.scala 80:57]
  wire [6:0] _sb_wmask_T_11 = 3'h6 == addr_low ? 7'h40 : {{1'd0}, _sb_wmask_T_9}; // @[Mux.scala 80:57]
  wire [7:0] sb_wmask = 3'h7 == addr_low ? 8'h80 : {{1'd0}, _sb_wmask_T_11}; // @[Mux.scala 80:57]
  wire [1:0] _sh_wmask_T_1 = 3'h0 == addr_low ? 2'h3 : 2'h0; // @[Mux.scala 80:57]
  wire [3:0] _sh_wmask_T_3 = 3'h2 == addr_low ? 4'hc : {{2'd0}, _sh_wmask_T_1}; // @[Mux.scala 80:57]
  wire [5:0] _sh_wmask_T_5 = 3'h4 == addr_low ? 6'h30 : {{2'd0}, _sh_wmask_T_3}; // @[Mux.scala 80:57]
  wire [7:0] sh_wmask = 3'h6 == addr_low ? 8'hc0 : {{2'd0}, _sh_wmask_T_5}; // @[Mux.scala 80:57]
  wire [3:0] _sw_wmask_T_1 = 3'h0 == addr_low ? 4'hf : 4'h0; // @[Mux.scala 80:57]
  wire [7:0] sw_wmask = 3'h4 == addr_low ? 8'hf0 : {{4'd0}, _sw_wmask_T_1}; // @[Mux.scala 80:57]
  wire [7:0] _dmem_wmask_T_1 = 4'h6 == io_lsu_op ? sb_wmask : 8'h0; // @[Mux.scala 80:57]
  wire [7:0] _dmem_wmask_T_3 = 4'h7 == io_lsu_op ? sh_wmask : _dmem_wmask_T_1; // @[Mux.scala 80:57]
  wire [7:0] _dmem_wmask_T_5 = 4'h8 == io_lsu_op ? sw_wmask : _dmem_wmask_T_3; // @[Mux.scala 80:57]
  wire [55:0] lb_rdata_hi = io_dmem_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo = io_dmem_rdata[7:0]; // @[LSU.scala 93:51]
  wire [63:0] _lb_rdata_T_2 = {lb_rdata_hi,lb_rdata_lo}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_1 = io_dmem_rdata[15] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_1 = io_dmem_rdata[15:8]; // @[LSU.scala 94:52]
  wire [63:0] _lb_rdata_T_5 = {lb_rdata_hi_1,lb_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_2 = io_dmem_rdata[23] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_2 = io_dmem_rdata[23:16]; // @[LSU.scala 95:52]
  wire [63:0] _lb_rdata_T_8 = {lb_rdata_hi_2,lb_rdata_lo_2}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_3 = io_dmem_rdata[31] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_3 = io_dmem_rdata[31:24]; // @[LSU.scala 96:52]
  wire [63:0] _lb_rdata_T_11 = {lb_rdata_hi_3,lb_rdata_lo_3}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_4 = io_dmem_rdata[39] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_4 = io_dmem_rdata[39:32]; // @[LSU.scala 97:52]
  wire [63:0] _lb_rdata_T_14 = {lb_rdata_hi_4,lb_rdata_lo_4}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_5 = io_dmem_rdata[47] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_5 = io_dmem_rdata[47:40]; // @[LSU.scala 98:52]
  wire [63:0] _lb_rdata_T_17 = {lb_rdata_hi_5,lb_rdata_lo_5}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_6 = io_dmem_rdata[55] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_6 = io_dmem_rdata[55:48]; // @[LSU.scala 99:52]
  wire [63:0] _lb_rdata_T_20 = {lb_rdata_hi_6,lb_rdata_lo_6}; // @[Cat.scala 30:58]
  wire [55:0] lb_rdata_hi_7 = io_dmem_rdata[63] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [7:0] lb_rdata_lo_7 = io_dmem_rdata[63:56]; // @[LSU.scala 100:52]
  wire [63:0] _lb_rdata_T_23 = {lb_rdata_hi_7,lb_rdata_lo_7}; // @[Cat.scala 30:58]
  wire [63:0] _lb_rdata_T_25 = 3'h1 == addr_low ? _lb_rdata_T_5 : _lb_rdata_T_2; // @[Mux.scala 80:57]
  wire [63:0] _lb_rdata_T_27 = 3'h2 == addr_low ? _lb_rdata_T_8 : _lb_rdata_T_25; // @[Mux.scala 80:57]
  wire [63:0] _lb_rdata_T_29 = 3'h3 == addr_low ? _lb_rdata_T_11 : _lb_rdata_T_27; // @[Mux.scala 80:57]
  wire [63:0] _lb_rdata_T_31 = 3'h4 == addr_low ? _lb_rdata_T_14 : _lb_rdata_T_29; // @[Mux.scala 80:57]
  wire [63:0] _lb_rdata_T_33 = 3'h5 == addr_low ? _lb_rdata_T_17 : _lb_rdata_T_31; // @[Mux.scala 80:57]
  wire [63:0] _lb_rdata_T_35 = 3'h6 == addr_low ? _lb_rdata_T_20 : _lb_rdata_T_33; // @[Mux.scala 80:57]
  wire [63:0] lb_rdata = 3'h7 == addr_low ? _lb_rdata_T_23 : _lb_rdata_T_35; // @[Mux.scala 80:57]
  wire [63:0] _lbu_rdata_T = {56'h0,lb_rdata_lo}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_1 = {56'h0,lb_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_2 = {56'h0,lb_rdata_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_3 = {56'h0,lb_rdata_lo_3}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_4 = {56'h0,lb_rdata_lo_4}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_5 = {56'h0,lb_rdata_lo_5}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_6 = {56'h0,lb_rdata_lo_6}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_7 = {56'h0,lb_rdata_lo_7}; // @[Cat.scala 30:58]
  wire [63:0] _lbu_rdata_T_9 = 3'h1 == addr_low ? _lbu_rdata_T_1 : _lbu_rdata_T; // @[Mux.scala 80:57]
  wire [63:0] _lbu_rdata_T_11 = 3'h2 == addr_low ? _lbu_rdata_T_2 : _lbu_rdata_T_9; // @[Mux.scala 80:57]
  wire [63:0] _lbu_rdata_T_13 = 3'h3 == addr_low ? _lbu_rdata_T_3 : _lbu_rdata_T_11; // @[Mux.scala 80:57]
  wire [63:0] _lbu_rdata_T_15 = 3'h4 == addr_low ? _lbu_rdata_T_4 : _lbu_rdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] _lbu_rdata_T_17 = 3'h5 == addr_low ? _lbu_rdata_T_5 : _lbu_rdata_T_15; // @[Mux.scala 80:57]
  wire [63:0] _lbu_rdata_T_19 = 3'h6 == addr_low ? _lbu_rdata_T_6 : _lbu_rdata_T_17; // @[Mux.scala 80:57]
  wire [63:0] lbu_rdata = 3'h7 == addr_low ? _lbu_rdata_T_7 : _lbu_rdata_T_19; // @[Mux.scala 80:57]
  wire [47:0] lh_rdata_hi = io_dmem_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] lh_rdata_lo = io_dmem_rdata[15:0]; // @[LSU.scala 114:52]
  wire [63:0] _lh_rdata_T_2 = {lh_rdata_hi,lh_rdata_lo}; // @[Cat.scala 30:58]
  wire [47:0] lh_rdata_hi_1 = io_dmem_rdata[31] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] lh_rdata_lo_1 = io_dmem_rdata[31:16]; // @[LSU.scala 115:52]
  wire [63:0] _lh_rdata_T_5 = {lh_rdata_hi_1,lh_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [47:0] lh_rdata_hi_2 = io_dmem_rdata[47] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] lh_rdata_lo_2 = io_dmem_rdata[47:32]; // @[LSU.scala 116:52]
  wire [63:0] _lh_rdata_T_8 = {lh_rdata_hi_2,lh_rdata_lo_2}; // @[Cat.scala 30:58]
  wire [47:0] lh_rdata_hi_3 = io_dmem_rdata[63] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [15:0] lh_rdata_lo_3 = io_dmem_rdata[63:48]; // @[LSU.scala 117:52]
  wire [63:0] _lh_rdata_T_11 = {lh_rdata_hi_3,lh_rdata_lo_3}; // @[Cat.scala 30:58]
  wire [63:0] _lh_rdata_T_13 = 3'h0 == addr_low ? _lh_rdata_T_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _lh_rdata_T_15 = 3'h2 == addr_low ? _lh_rdata_T_5 : _lh_rdata_T_13; // @[Mux.scala 80:57]
  wire [63:0] _lh_rdata_T_17 = 3'h4 == addr_low ? _lh_rdata_T_8 : _lh_rdata_T_15; // @[Mux.scala 80:57]
  wire [63:0] lh_rdata = 3'h6 == addr_low ? _lh_rdata_T_11 : _lh_rdata_T_17; // @[Mux.scala 80:57]
  wire [63:0] _lhu_rdata_T = {48'h0,lh_rdata_lo}; // @[Cat.scala 30:58]
  wire [63:0] _lhu_rdata_T_1 = {48'h0,lh_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _lhu_rdata_T_2 = {48'h0,lh_rdata_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _lhu_rdata_T_3 = {48'h0,lh_rdata_lo_3}; // @[Cat.scala 30:58]
  wire [63:0] _lhu_rdata_T_5 = 3'h0 == addr_low ? _lhu_rdata_T : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _lhu_rdata_T_7 = 3'h2 == addr_low ? _lhu_rdata_T_1 : _lhu_rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _lhu_rdata_T_9 = 3'h4 == addr_low ? _lhu_rdata_T_2 : _lhu_rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] lhu_rdata = 3'h6 == addr_low ? _lhu_rdata_T_3 : _lhu_rdata_T_9; // @[Mux.scala 80:57]
  wire [31:0] lw_rdata_hi = io_dmem_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] lw_rdata_lo = io_dmem_rdata[31:0]; // @[LSU.scala 126:52]
  wire [63:0] _lw_rdata_T_2 = {lw_rdata_hi,lw_rdata_lo}; // @[Cat.scala 30:58]
  wire [31:0] lw_rdata_hi_1 = io_dmem_rdata[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] lw_rdata_lo_1 = io_dmem_rdata[63:32]; // @[LSU.scala 127:52]
  wire [63:0] _lw_rdata_T_5 = {lw_rdata_hi_1,lw_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _lw_rdata_T_7 = 3'h0 == addr_low ? _lw_rdata_T_2 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] lw_rdata = 3'h4 == addr_low ? _lw_rdata_T_5 : _lw_rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _lwu_rdata_T = {32'h0,lw_rdata_lo}; // @[Cat.scala 30:58]
  wire [63:0] _lwu_rdata_T_1 = {32'h0,lw_rdata_lo_1}; // @[Cat.scala 30:58]
  wire [63:0] _lwu_rdata_T_3 = 3'h0 == addr_low ? _lwu_rdata_T : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] lwu_rdata = 3'h4 == addr_low ? _lwu_rdata_T_1 : _lwu_rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _load_rdata_T_1 = 4'h1 == io_lsu_op ? lb_rdata : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _load_rdata_T_3 = 4'h4 == io_lsu_op ? lbu_rdata : _load_rdata_T_1; // @[Mux.scala 80:57]
  wire [63:0] _load_rdata_T_5 = 4'h2 == io_lsu_op ? lh_rdata : _load_rdata_T_3; // @[Mux.scala 80:57]
  wire [63:0] _load_rdata_T_7 = 4'h5 == io_lsu_op ? lhu_rdata : _load_rdata_T_5; // @[Mux.scala 80:57]
  wire [63:0] _load_rdata_T_9 = 4'h3 == io_lsu_op ? lw_rdata : _load_rdata_T_7; // @[Mux.scala 80:57]
  wire [63:0] _load_rdata_T_11 = 4'h9 == io_lsu_op ? lwu_rdata : _load_rdata_T_9; // @[Mux.scala 80:57]
  reg [2:0] state; // @[LSU.scala 155:22]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_0 = io_is_lsu ? 3'h3 : 3'h0; // @[LSU.scala 168:28 LSU.scala 169:15 LSU.scala 172:15]
  wire  _GEN_3 = io_is_lsu & io_is_mdu | io_is_lsu; // @[LSU.scala 165:38 LSU.scala 167:23]
  wire  _GEN_5 = fence_i ? 1'h0 : _GEN_3; // @[LSU.scala 162:20 LSU.scala 164:23]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_6 = io_dmem_data_ok ? 3'h2 : state; // @[LSU.scala 184:37 LSU.scala 185:15 LSU.scala 155:22]
  wire  _GEN_7 = io_dmem_data_ok ? 1'h0 : 1'h1; // @[LSU.scala 184:37 LSU.scala 186:23 LSU.scala 177:21]
  wire [2:0] _GEN_8 = io_mdu_ok ? 3'h3 : _GEN_6; // @[LSU.scala 181:28 LSU.scala 182:15]
  wire  _GEN_9 = io_mdu_ok | _GEN_7; // @[LSU.scala 181:28 LSU.scala 183:23]
  wire  _GEN_11 = io_dmem_data_ok & io_mdu_ok ? 1'h0 : _GEN_9; // @[LSU.scala 178:40 LSU.scala 180:23]
  wire  _T_4 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_12 = io_dmem_data_ok ? 3'h0 : state; // @[LSU.scala 191:30 LSU.scala 192:15 LSU.scala 155:22]
  wire  _T_5 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_13 = io_mdu_ok ? 3'h0 : state; // @[LSU.scala 198:21 LSU.scala 199:15 LSU.scala 155:22]
  wire  _T_6 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  dcache_fence_finish = io_dmem_fence_finish; // @[LSU.scala 150:33 LSU.scala 151:23]
  wire [2:0] _GEN_14 = icache_fence_finish_0 ? 3'h6 : state; // @[LSU.scala 210:41 LSU.scala 211:15 LSU.scala 155:22]
  wire  _GEN_15 = dcache_fence_finish ? 1'h0 : 1'h1; // @[LSU.scala 207:41 LSU.scala 208:23 LSU.scala 203:21]
  wire [2:0] _GEN_16 = dcache_fence_finish ? 3'h5 : _GEN_14; // @[LSU.scala 207:41 LSU.scala 209:15]
  wire  _GEN_17 = dcache_fence_finish & icache_fence_finish_0 ? 1'h0 : _GEN_15; // @[LSU.scala 204:57 LSU.scala 205:23]
  wire [2:0] _GEN_18 = dcache_fence_finish & icache_fence_finish_0 ? 3'h0 : _GEN_16; // @[LSU.scala 204:57 LSU.scala 206:15]
  wire  _T_8 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_19 = icache_fence_finish_0 ? 3'h0 : state; // @[LSU.scala 215:34 LSU.scala 216:15 LSU.scala 155:22]
  wire  _T_9 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_21 = _T_9 ? 3'h0 : state; // @[Conditional.scala 39:67 LSU.scala 221:13 LSU.scala 155:22]
  wire [2:0] _GEN_22 = _T_8 ? _GEN_19 : _GEN_21; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_25 = _T_6 ? _GEN_18 : _GEN_22; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_27 = _T_5 ? _GEN_13 : _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_28 = _T_5 ? 1'h0 : _T_6 & _GEN_17; // @[Conditional.scala 39:67 LSU.scala 158:17]
  wire  _GEN_31 = _T_4 ? 1'h0 : _GEN_28; // @[Conditional.scala 39:67 LSU.scala 158:17]
  wire  _GEN_32 = _T_2 ? _GEN_11 : _T_4 & _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_2 ? 1'h0 : _GEN_31; // @[Conditional.scala 39:67 LSU.scala 158:17]
  assign io_dmem_valid = _T ? _GEN_5 : _GEN_32; // @[Conditional.scala 40:58]
  assign io_dmem_op = io_wen ? 1'h0 : 1'h1; // @[LSU.scala 225:20]
  assign io_dmem_addr = io_addr; // @[LSU.scala 226:16]
  assign io_dmem_wstrb = 4'hb == io_lsu_op ? 8'hff : _dmem_wmask_T_5; // @[Mux.scala 80:57]
  assign io_dmem_wdata = 4'hb == io_lsu_op ? io_wdata : _dmem_wdata_T_5; // @[Mux.scala 80:57]
  assign io_dmem_fence = _T ? 1'h0 : _GEN_34; // @[Conditional.scala 40:58 LSU.scala 158:17]
  assign io_addr = _io_addr_T_1[31:0]; // @[LSU.scala 28:33]
  assign io_rdata = 4'ha == io_lsu_op ? io_dmem_rdata : _load_rdata_T_11; // @[Mux.scala 80:57]
  assign dcache_fence_finish_0 = dcache_fence_finish;
  always @(posedge clock) begin
    if (reset) begin // @[LSU.scala 155:22]
      state <= 3'h0; // @[LSU.scala 155:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (fence_i) begin // @[LSU.scala 162:20]
        state <= 3'h4; // @[LSU.scala 163:15]
      end else if (io_is_lsu & io_is_mdu) begin // @[LSU.scala 165:38]
        state <= 3'h1; // @[LSU.scala 166:15]
      end else begin
        state <= _GEN_0;
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (io_dmem_data_ok & io_mdu_ok) begin // @[LSU.scala 178:40]
        state <= 3'h0; // @[LSU.scala 179:15]
      end else begin
        state <= _GEN_8;
      end
    end else if (_T_4) begin // @[Conditional.scala 39:67]
      state <= _GEN_12;
    end else begin
      state <= _GEN_27;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         reset,
  input  [31:0] io_pc,
  input  [2:0]  io_csr_op,
  input  [11:0] io_addr,
  input  [63:0] io_src,
  output [63:0] io_rdata,
  output        io_is_reflush,
  output [31:0] io_csr_target,
  output        io_handle_int,
  input         io_valid,
  input         clint_has_int
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mcycle; // @[CSR.scala 28:23]
  reg [63:0] mepc; // @[CSR.scala 29:21]
  reg [63:0] mcause; // @[CSR.scala 30:23]
  reg [63:0] mstatus; // @[CSR.scala 31:24]
  reg [63:0] mtvec; // @[CSR.scala 32:22]
  reg [63:0] mip; // @[CSR.scala 33:20]
  reg [63:0] mie; // @[CSR.scala 34:20]
  reg [63:0] mscratch; // @[CSR.scala 35:25]
  wire  wen = io_csr_op == 3'h1 | io_csr_op == 3'h2 | io_csr_op == 3'h3; // @[CSR.scala 43:59]
  wire  _T_36 = io_addr == 12'h342; // @[MAP.scala 23:18]
  wire  _T_33 = io_addr == 12'h340; // @[MAP.scala 23:18]
  wire  _T_30 = io_addr == 12'hb00; // @[MAP.scala 23:18]
  wire  _T_27 = io_addr == 12'h304; // @[MAP.scala 23:18]
  wire  _T_24 = io_addr == 12'h344; // @[MAP.scala 23:18]
  wire  _T_21 = io_addr == 12'h300; // @[MAP.scala 23:18]
  wire  _T_18 = io_addr == 12'h305; // @[MAP.scala 23:18]
  wire  _T_15 = io_addr == 12'h341; // @[MAP.scala 23:18]
  wire [63:0] _GEN_14 = io_addr == 12'h341 ? mepc : 64'h0; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _GEN_16 = io_addr == 12'h305 ? mtvec : _GEN_14; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _GEN_18 = io_addr == 12'h300 ? mstatus : _GEN_16; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _GEN_20 = io_addr == 12'h344 ? mip : _GEN_18; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _GEN_22 = io_addr == 12'h304 ? mie : _GEN_20; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _GEN_24 = io_addr == 12'hb00 ? mcycle : _GEN_22; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _GEN_26 = io_addr == 12'h340 ? mscratch : _GEN_24; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] rdata = io_addr == 12'h342 ? mcause : _GEN_26; // @[MAP.scala 23:25 MAP.scala 24:15]
  wire [63:0] _wdata_T = rdata | io_src; // @[CSR.scala 63:25]
  wire [63:0] _wdata_T_1 = ~io_src; // @[CSR.scala 64:28]
  wire [63:0] _wdata_T_2 = rdata & _wdata_T_1; // @[CSR.scala 64:25]
  wire [63:0] _wdata_T_4 = 3'h1 == io_csr_op ? io_src : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _wdata_T_6 = 3'h2 == io_csr_op ? _wdata_T : _wdata_T_4; // @[Mux.scala 80:57]
  wire [63:0] wdata = 3'h3 == io_csr_op ? _wdata_T_2 : _wdata_T_6; // @[Mux.scala 80:57]
  wire  _T_13 = io_csr_op == 3'h4; // @[CSR.scala 67:16]
  wire [55:0] mstatus_hi_hi_hi = mstatus[63:8]; // @[CSR.scala 70:27]
  wire  mstatus_hi_hi_lo = mstatus[3]; // @[CSR.scala 70:43]
  wire [2:0] mstatus_hi_lo = mstatus[6:4]; // @[CSR.scala 70:55]
  wire [2:0] mstatus_lo_lo = mstatus[2:0]; // @[CSR.scala 70:75]
  wire [63:0] _mstatus_T = {mstatus_hi_hi_hi,mstatus_hi_hi_lo,mstatus_hi_lo,1'h0,mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [29:0] csr_target_hi = mtvec[31:2]; // @[CSR.scala 72:28]
  wire [31:0] _csr_target_T = {csr_target_hi,2'h0}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_2 = io_csr_op == 3'h4 ? _mstatus_T : mstatus; // @[CSR.scala 67:31 CSR.scala 70:13 CSR.scala 31:24]
  wire [31:0] _GEN_4 = io_csr_op == 3'h4 ? _csr_target_T : 32'h0; // @[CSR.scala 67:31 CSR.scala 72:16]
  wire  handle_int = clint_has_int & mstatus_hi_hi_lo & mie[7] & io_valid; // @[CSR.scala 96:40]
  wire  _GEN_9 = handle_int | _T_13; // @[CSR.scala 75:20 CSR.scala 80:15]
  wire [31:0] _GEN_10 = handle_int ? _csr_target_T : _GEN_4; // @[CSR.scala 75:20 CSR.scala 81:16]
  wire  mstatus_lo_hi = mstatus[7]; // @[CSR.scala 85:63]
  wire [63:0] _mstatus_T_2 = {mstatus_hi_hi_hi,1'h1,mstatus_hi_lo,mstatus_lo_hi,mstatus_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mcycle_T_1 = mcycle + 64'h1; // @[CSR.scala 90:20]
  wire [63:0] _mepc_T = wdata & 64'hfffffffffffffffc; // @[MAP.scala 10:14]
  wire [63:0] _mepc_T_2 = mepc & 64'h3; // @[MAP.scala 10:33]
  wire [63:0] _mepc_T_3 = _mepc_T | _mepc_T_2; // @[MAP.scala 10:22]
  wire  mstatus_mstatus_new_hi = wdata[16:15] == 2'h3 | wdata[14:13] == 2'h3; // @[CSR.scala 46:57]
  wire [62:0] mstatus_mstatus_new_lo = wdata[62:0]; // @[CSR.scala 46:98]
  wire [63:0] mstatus_mstatus_new = {mstatus_mstatus_new_hi,mstatus_mstatus_new_lo}; // @[Cat.scala 30:58]
  wire [63:0] _mip_T_2 = mip & 64'h1; // @[MAP.scala 10:33]
  wire [55:0] mip_hi_hi = mip[63:8]; // @[CSR.scala 98:19]
  wire [6:0] mip_lo = mip[6:0]; // @[CSR.scala 98:36]
  wire [63:0] _mip_T_4 = {mip_hi_hi,1'h1,mip_lo}; // @[Cat.scala 30:58]
  assign io_rdata = io_addr == 12'h342 ? mcause : _GEN_26; // @[MAP.scala 23:25 MAP.scala 24:15]
  assign io_is_reflush = io_csr_op == 3'h5 | _GEN_9; // @[CSR.scala 84:30 CSR.scala 86:15]
  assign io_csr_target = io_csr_op == 3'h5 ? mepc[31:0] : _GEN_10; // @[CSR.scala 84:30 CSR.scala 87:16]
  assign io_handle_int = clint_has_int & mstatus_hi_hi_lo & mie[7] & io_valid; // @[CSR.scala 96:40]
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 28:23]
      mcycle <= 64'h0; // @[CSR.scala 28:23]
    end else if (_T_30 & wen) begin // @[MAP.scala 27:34]
      if (3'h3 == io_csr_op) begin // @[Mux.scala 80:57]
        mcycle <= _wdata_T_2;
      end else if (3'h2 == io_csr_op) begin // @[Mux.scala 80:57]
        mcycle <= _wdata_T;
      end else begin
        mcycle <= _wdata_T_4;
      end
    end else begin
      mcycle <= _mcycle_T_1; // @[CSR.scala 90:10]
    end
    if (reset) begin // @[CSR.scala 29:21]
      mepc <= 64'h0; // @[CSR.scala 29:21]
    end else if (_T_15 & wen) begin // @[MAP.scala 27:34]
      mepc <= _mepc_T_3; // @[MAP.scala 28:13]
    end else if (handle_int) begin // @[CSR.scala 75:20]
      mepc <= {{32'd0}, io_pc}; // @[CSR.scala 77:10]
    end else if (io_csr_op == 3'h4) begin // @[CSR.scala 67:31]
      mepc <= {{32'd0}, io_pc}; // @[CSR.scala 68:10]
    end
    if (reset) begin // @[CSR.scala 30:23]
      mcause <= 64'h0; // @[CSR.scala 30:23]
    end else if (_T_36 & wen) begin // @[MAP.scala 27:34]
      if (3'h3 == io_csr_op) begin // @[Mux.scala 80:57]
        mcause <= _wdata_T_2;
      end else if (3'h2 == io_csr_op) begin // @[Mux.scala 80:57]
        mcause <= _wdata_T;
      end else begin
        mcause <= _wdata_T_4;
      end
    end else if (handle_int) begin // @[CSR.scala 75:20]
      mcause <= 64'h8000000000000007; // @[CSR.scala 78:12]
    end else if (io_csr_op == 3'h4) begin // @[CSR.scala 67:31]
      mcause <= 64'hb; // @[CSR.scala 69:12]
    end
    if (reset) begin // @[CSR.scala 31:24]
      mstatus <= 64'h1800; // @[CSR.scala 31:24]
    end else if (_T_21 & wen) begin // @[MAP.scala 27:34]
      mstatus <= mstatus_mstatus_new; // @[MAP.scala 28:13]
    end else if (io_csr_op == 3'h5) begin // @[CSR.scala 84:30]
      mstatus <= _mstatus_T_2; // @[CSR.scala 85:13]
    end else if (handle_int) begin // @[CSR.scala 75:20]
      mstatus <= _mstatus_T; // @[CSR.scala 79:13]
    end else begin
      mstatus <= _GEN_2;
    end
    if (reset) begin // @[CSR.scala 32:22]
      mtvec <= 64'h0; // @[CSR.scala 32:22]
    end else if (_T_18 & wen) begin // @[MAP.scala 27:34]
      if (3'h3 == io_csr_op) begin // @[Mux.scala 80:57]
        mtvec <= _wdata_T_2;
      end else if (3'h2 == io_csr_op) begin // @[Mux.scala 80:57]
        mtvec <= _wdata_T;
      end else begin
        mtvec <= _wdata_T_4;
      end
    end
    if (reset) begin // @[CSR.scala 33:20]
      mip <= 64'h0; // @[CSR.scala 33:20]
    end else if (handle_int) begin // @[CSR.scala 96:53]
      mip <= _mip_T_4; // @[CSR.scala 98:9]
    end else if (_T_24 & wen) begin // @[MAP.scala 27:34]
      mip <= _mip_T_2; // @[MAP.scala 28:13]
    end else if (handle_int) begin // @[CSR.scala 75:20]
      mip <= 64'h0; // @[CSR.scala 76:9]
    end
    if (reset) begin // @[CSR.scala 34:20]
      mie <= 64'h0; // @[CSR.scala 34:20]
    end else if (_T_27 & wen) begin // @[MAP.scala 27:34]
      if (3'h3 == io_csr_op) begin // @[Mux.scala 80:57]
        mie <= _wdata_T_2;
      end else if (3'h2 == io_csr_op) begin // @[Mux.scala 80:57]
        mie <= _wdata_T;
      end else begin
        mie <= _wdata_T_4;
      end
    end
    if (reset) begin // @[CSR.scala 35:25]
      mscratch <= 64'h0; // @[CSR.scala 35:25]
    end else if (_T_33 & wen) begin // @[MAP.scala 27:34]
      if (3'h3 == io_csr_op) begin // @[Mux.scala 80:57]
        mscratch <= _wdata_T_2;
      end else if (3'h2 == io_csr_op) begin // @[Mux.scala 80:57]
        mscratch <= _wdata_T;
      end else begin
        mscratch <= _wdata_T_4;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mcycle = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mepc = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mstatus = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mtvec = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mip = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mie = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  mscratch = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLINT(
  input         clock,
  input         reset,
  input         io_is_mtime,
  input         io_is_mtimecmp,
  input         io_is_clint,
  input         io_wen,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output        has_int_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[CLINT.scala 17:22]
  reg [63:0] mtimecmp; // @[CLINT.scala 18:25]
  reg  count_2; // @[CLINT.scala 27:24]
  wire [63:0] _mtime_T_1 = mtime + 64'h1; // @[CLINT.scala 31:20]
  wire [63:0] _GEN_0 = ~count_2 ? _mtime_T_1 : mtime; // @[CLINT.scala 30:26 CLINT.scala 31:11 CLINT.scala 17:22]
  wire [63:0] _rdata_T = io_is_mtime ? mtime : mtimecmp; // @[CLINT.scala 37:19]
  wire [63:0] _GEN_1 = io_wen ? _rdata_T : 64'h0; // @[CLINT.scala 36:16 CLINT.scala 37:13]
  wire  _GEN_9 = mtime >= mtimecmp; // @[CLINT.scala 51:15]
  wire  has_int = mtime >= mtimecmp; // @[CLINT.scala 51:15]
  assign io_rdata = io_is_clint ? _GEN_1 : 64'h0; // @[CLINT.scala 35:19]
  assign has_int_0 = _GEN_9;
  always @(posedge clock) begin
    if (reset) begin // @[CLINT.scala 17:22]
      mtime <= 64'h0; // @[CLINT.scala 17:22]
    end else if (io_is_clint) begin // @[CLINT.scala 35:19]
      if (~io_wen) begin // @[CLINT.scala 39:17]
        if (io_is_mtime) begin // @[CLINT.scala 40:23]
          mtime <= io_wdata; // @[CLINT.scala 41:15]
        end else begin
          mtime <= _GEN_0;
        end
      end else begin
        mtime <= _GEN_0;
      end
    end else begin
      mtime <= _GEN_0;
    end
    if (reset) begin // @[CLINT.scala 18:25]
      mtimecmp <= 64'h0; // @[CLINT.scala 18:25]
    end else if (io_is_clint) begin // @[CLINT.scala 35:19]
      if (~io_wen) begin // @[CLINT.scala 39:17]
        if (io_is_mtimecmp) begin // @[CLINT.scala 43:26]
          mtimecmp <= io_wdata; // @[CLINT.scala 44:18]
        end
      end
    end
    if (reset) begin // @[CLINT.scala 27:24]
      count_2 <= 1'h0; // @[CLINT.scala 27:24]
    end else begin
      count_2 <= count_2 + 1'h1; // @[CLINT.scala 28:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  count_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io_dmem_valid,
  output        io_dmem_op,
  output [31:0] io_dmem_addr,
  output [7:0]  io_dmem_wstrb,
  output [63:0] io_dmem_wdata,
  output        io_dmem_fence,
  input         io_dmem_fence_finish,
  input         io_dmem_data_ok,
  input  [63:0] io_dmem_rdata,
  output        io_in_ready,
  input         io_in_valid,
  input         io_in_bits_0_valid,
  input  [31:0] io_in_bits_0_pc,
  input  [31:0] io_in_bits_0_inst,
  input  [63:0] io_in_bits_0_src1_value,
  input  [63:0] io_in_bits_0_src2_value,
  input  [63:0] io_in_bits_0_rs2_value,
  input  [63:0] io_in_bits_0_imm,
  input  [4:0]  io_in_bits_0_rs1,
  input  [4:0]  io_in_bits_0_dest,
  input  [2:0]  io_in_bits_0_fu_type,
  input  [3:0]  io_in_bits_0_bru_op,
  input  [4:0]  io_in_bits_0_alu_op,
  input  [3:0]  io_in_bits_0_lsu_op,
  input  [2:0]  io_in_bits_0_csr_op,
  input  [3:0]  io_in_bits_0_mdu_op,
  input         io_in_bits_0_wen,
  input         io_in_bits_0_rv64,
  input         io_in_bits_0_bp_br_taken,
  input  [31:0] io_in_bits_0_bp_br_target,
  input  [1:0]  io_in_bits_0_bp_br_type,
  input         io_in_bits_1_valid,
  input  [31:0] io_in_bits_1_pc,
  input  [31:0] io_in_bits_1_inst,
  input  [63:0] io_in_bits_1_src1_value,
  input  [63:0] io_in_bits_1_src2_value,
  input  [63:0] io_in_bits_1_rs2_value,
  input  [63:0] io_in_bits_1_imm,
  input  [4:0]  io_in_bits_1_rs1,
  input  [4:0]  io_in_bits_1_dest,
  input  [2:0]  io_in_bits_1_fu_type,
  input  [3:0]  io_in_bits_1_bru_op,
  input  [4:0]  io_in_bits_1_alu_op,
  input  [3:0]  io_in_bits_1_lsu_op,
  input  [2:0]  io_in_bits_1_csr_op,
  input  [3:0]  io_in_bits_1_mdu_op,
  input         io_in_bits_1_wen,
  input         io_in_bits_1_rv64,
  input         io_in_bits_1_bp_br_taken,
  input  [31:0] io_in_bits_1_bp_br_target,
  input  [1:0]  io_in_bits_1_bp_br_type,
  output        io_out_valid,
  output        io_out_bits_0_valid,
  output [31:0] io_out_bits_0_pc,
  output [63:0] io_out_bits_0_final_result,
  output [4:0]  io_out_bits_0_dest,
  output        io_out_bits_0_wen,
  output        io_out_bits_1_valid,
  output [63:0] io_out_bits_1_final_result,
  output [4:0]  io_out_bits_1_dest,
  output        io_out_bits_1_wen,
  output        io_forward_0_blk_valid,
  output        io_forward_0_fwd_valid,
  output [4:0]  io_forward_0_rf_waddr,
  output [63:0] io_forward_0_rf_wdata,
  output        io_forward_1_blk_valid,
  output        io_forward_1_fwd_valid,
  output [4:0]  io_forward_1_rf_waddr,
  output [63:0] io_forward_1_rf_wdata,
  output        io_reflush_bus_is_reflush,
  output [31:0] io_reflush_bus_br_target,
  output        io_bpu_valid,
  output [31:0] io_bpu_pc,
  output        io_bpu_bp_taken,
  output [31:0] io_bpu_bp_target,
  output [1:0]  io_bpu_bp_type,
  output        io_bpu_bp_wrong,
  output        io_bpu_fence,
  output [2:0]  io_bpu_call_count,
  output [2:0]  io_bpu_ret_count,
  output        frontend_reflush_0,
  output        dcache_fence_finish,
  output        fence_0,
  input         icache_fence_finish
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] alu_0_io_alu_op; // @[EXU.scala 20:21]
  wire  alu_0_io_rv64; // @[EXU.scala 20:21]
  wire [63:0] alu_0_io_src1; // @[EXU.scala 20:21]
  wire [63:0] alu_0_io_src2; // @[EXU.scala 20:21]
  wire [63:0] alu_0_io_result; // @[EXU.scala 20:21]
  wire [4:0] alu_1_io_alu_op; // @[EXU.scala 20:21]
  wire  alu_1_io_rv64; // @[EXU.scala 20:21]
  wire [63:0] alu_1_io_src1; // @[EXU.scala 20:21]
  wire [63:0] alu_1_io_src2; // @[EXU.scala 20:21]
  wire [63:0] alu_1_io_result; // @[EXU.scala 20:21]
  wire  mdu_clock; // @[EXU.scala 23:19]
  wire  mdu_reset; // @[EXU.scala 23:19]
  wire [3:0] mdu_io_mdu_op; // @[EXU.scala 23:19]
  wire  mdu_io_rv64; // @[EXU.scala 23:19]
  wire [63:0] mdu_io_src1; // @[EXU.scala 23:19]
  wire [63:0] mdu_io_src2; // @[EXU.scala 23:19]
  wire  mdu_io_result_ok; // @[EXU.scala 23:19]
  wire [63:0] mdu_io_result; // @[EXU.scala 23:19]
  wire [3:0] bru_io_bru_op; // @[EXU.scala 24:19]
  wire [63:0] bru_io_src1; // @[EXU.scala 24:19]
  wire [63:0] bru_io_src2; // @[EXU.scala 24:19]
  wire [31:0] bru_io_pc; // @[EXU.scala 24:19]
  wire [63:0] bru_io_imm; // @[EXU.scala 24:19]
  wire  bru_io_br_taken; // @[EXU.scala 24:19]
  wire [31:0] bru_io_br_target; // @[EXU.scala 24:19]
  wire [4:0] bru_io_rs1; // @[EXU.scala 24:19]
  wire [4:0] bru_io_rd; // @[EXU.scala 24:19]
  wire [1:0] bru_io_btb_type; // @[EXU.scala 24:19]
  wire  lsu_clock; // @[EXU.scala 25:19]
  wire  lsu_reset; // @[EXU.scala 25:19]
  wire  lsu_io_dmem_valid; // @[EXU.scala 25:19]
  wire  lsu_io_dmem_op; // @[EXU.scala 25:19]
  wire [31:0] lsu_io_dmem_addr; // @[EXU.scala 25:19]
  wire [7:0] lsu_io_dmem_wstrb; // @[EXU.scala 25:19]
  wire [63:0] lsu_io_dmem_wdata; // @[EXU.scala 25:19]
  wire  lsu_io_dmem_fence; // @[EXU.scala 25:19]
  wire  lsu_io_dmem_fence_finish; // @[EXU.scala 25:19]
  wire  lsu_io_dmem_data_ok; // @[EXU.scala 25:19]
  wire [63:0] lsu_io_dmem_rdata; // @[EXU.scala 25:19]
  wire [63:0] lsu_io_src1; // @[EXU.scala 25:19]
  wire [63:0] lsu_io_src2; // @[EXU.scala 25:19]
  wire [63:0] lsu_io_wdata; // @[EXU.scala 25:19]
  wire [31:0] lsu_io_addr; // @[EXU.scala 25:19]
  wire  lsu_io_is_lsu; // @[EXU.scala 25:19]
  wire  lsu_io_wen; // @[EXU.scala 25:19]
  wire [3:0] lsu_io_lsu_op; // @[EXU.scala 25:19]
  wire [63:0] lsu_io_rdata; // @[EXU.scala 25:19]
  wire  lsu_io_is_mdu; // @[EXU.scala 25:19]
  wire  lsu_io_mdu_ok; // @[EXU.scala 25:19]
  wire  lsu_dcache_fence_finish_0; // @[EXU.scala 25:19]
  wire  lsu_fence_i; // @[EXU.scala 25:19]
  wire  lsu_icache_fence_finish_0; // @[EXU.scala 25:19]
  wire  csr_clock; // @[EXU.scala 26:19]
  wire  csr_reset; // @[EXU.scala 26:19]
  wire [31:0] csr_io_pc; // @[EXU.scala 26:19]
  wire [2:0] csr_io_csr_op; // @[EXU.scala 26:19]
  wire [11:0] csr_io_addr; // @[EXU.scala 26:19]
  wire [63:0] csr_io_src; // @[EXU.scala 26:19]
  wire [63:0] csr_io_rdata; // @[EXU.scala 26:19]
  wire  csr_io_is_reflush; // @[EXU.scala 26:19]
  wire [31:0] csr_io_csr_target; // @[EXU.scala 26:19]
  wire  csr_io_handle_int; // @[EXU.scala 26:19]
  wire  csr_io_valid; // @[EXU.scala 26:19]
  wire  csr_clint_has_int; // @[EXU.scala 26:19]
  wire  clint_clock; // @[EXU.scala 27:21]
  wire  clint_reset; // @[EXU.scala 27:21]
  wire  clint_io_is_mtime; // @[EXU.scala 27:21]
  wire  clint_io_is_mtimecmp; // @[EXU.scala 27:21]
  wire  clint_io_is_clint; // @[EXU.scala 27:21]
  wire  clint_io_wen; // @[EXU.scala 27:21]
  wire [63:0] clint_io_wdata; // @[EXU.scala 27:21]
  wire [63:0] clint_io_rdata; // @[EXU.scala 27:21]
  wire  clint_has_int_0; // @[EXU.scala 27:21]
  reg [1:0] blk_state; // @[EXU.scala 51:26]
  wire  _GEN_0 = io_in_bits_0_fu_type == 3'h4 & io_in_bits_0_valid & io_in_valid; // @[EXU.scala 72:61 EXU.scala 73:14 EXU.scala 64:10]
  wire  is_mdu = io_in_bits_1_fu_type == 3'h4 & io_in_bits_1_valid ? io_in_valid : _GEN_0; // @[EXU.scala 72:61 EXU.scala 73:14]
  wire [3:0] _mdu_io_mdu_op_T_1 = is_mdu ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [3:0] _mdu_io_mdu_op_T_2 = io_in_bits_0_mdu_op & _mdu_io_mdu_op_T_1; // @[EXU.scala 76:42]
  wire [63:0] _GEN_1 = io_in_bits_0_fu_type == 3'h4 & io_in_bits_0_valid ? io_in_bits_0_src1_value : 64'h0; // @[EXU.scala 72:61 EXU.scala 74:19 EXU.scala 65:15]
  wire [63:0] _GEN_2 = io_in_bits_0_fu_type == 3'h4 & io_in_bits_0_valid ? io_in_bits_0_src2_value : 64'h0; // @[EXU.scala 72:61 EXU.scala 75:19 EXU.scala 66:15]
  wire [3:0] _GEN_3 = io_in_bits_0_fu_type == 3'h4 & io_in_bits_0_valid ? _mdu_io_mdu_op_T_2 : 4'h0; // @[EXU.scala 72:61 EXU.scala 76:21 EXU.scala 67:17]
  wire  _GEN_4 = io_in_bits_0_fu_type == 3'h4 & io_in_bits_0_valid & io_in_bits_0_rv64; // @[EXU.scala 72:61 EXU.scala 77:19 EXU.scala 68:15]
  wire [3:0] _mdu_io_mdu_op_T_5 = io_in_bits_1_mdu_op & _mdu_io_mdu_op_T_1; // @[EXU.scala 76:42]
  wire  _T_4 = io_in_bits_0_fu_type == 3'h1; // @[EXU.scala 94:30]
  wire  _T_5 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid; // @[EXU.scala 94:41]
  wire [3:0] _GEN_10 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_bru_op : 4'h0; // @[EXU.scala 94:62 EXU.scala 95:21 EXU.scala 86:17]
  wire [63:0] _GEN_11 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_src1_value : 64'h0; // @[EXU.scala 94:62 EXU.scala 96:19 EXU.scala 87:15]
  wire [63:0] _GEN_12 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_src2_value : 64'h0; // @[EXU.scala 94:62 EXU.scala 97:19 EXU.scala 88:15]
  wire [31:0] _GEN_13 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_pc : 32'h0; // @[EXU.scala 94:62 EXU.scala 98:17 EXU.scala 89:13]
  wire [63:0] _GEN_14 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_imm : 64'h0; // @[EXU.scala 94:62 EXU.scala 99:18 EXU.scala 90:14]
  wire [4:0] _GEN_15 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_rs1 : 5'h0; // @[EXU.scala 94:62 EXU.scala 100:18 EXU.scala 91:14]
  wire [4:0] _GEN_16 = io_in_bits_0_fu_type == 3'h1 & io_in_bits_0_valid ? io_in_bits_0_dest : 5'h0; // @[EXU.scala 94:62 EXU.scala 101:17 EXU.scala 92:13]
  wire  _T_6 = io_in_bits_1_fu_type == 3'h1; // @[EXU.scala 94:30]
  wire  _T_7 = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid; // @[EXU.scala 94:41]
  reg [2:0] call_count; // @[EXU.scala 106:27]
  reg [2:0] ret_count; // @[EXU.scala 107:26]
  wire [1:0] br_type = bru_io_btb_type; // @[EXU.scala 42:21 EXU.scala 84:11]
  wire [2:0] _GEN_106 = {{2'd0}, br_type == 2'h0}; // @[EXU.scala 113:30]
  wire [2:0] _call_count_T_2 = call_count + _GEN_106; // @[EXU.scala 113:30]
  wire [2:0] _GEN_107 = {{2'd0}, br_type == 2'h1}; // @[EXU.scala 114:28]
  wire [2:0] _ret_count_T_2 = ret_count + _GEN_107; // @[EXU.scala 114:28]
  wire  csr_is_reflush = csr_io_is_reflush; // @[EXU.scala 43:28 EXU.scala 171:18]
  wire  handle_int = csr_io_handle_int; // @[EXU.scala 45:24 EXU.scala 173:14]
  wire  _frontend_reflush_T = ~handle_int; // @[EXU.scala 228:44]
  wire  fence = csr_io_csr_op == 3'h6; // @[EXU.scala 174:27]
  wire  br_taken = bru_io_br_taken; // @[EXU.scala 40:22 EXU.scala 82:12]
  wire [31:0] br_target = bru_io_br_target; // @[EXU.scala 41:23 EXU.scala 83:13]
  wire  _bp_wrong_T_13 = br_taken & io_in_bits_1_bp_br_taken & (br_target != io_in_bits_1_bp_br_target | br_type !=
    io_in_bits_1_bp_br_type); // @[EXU.scala 132:45]
  wire  _bp_wrong_T_14 = br_taken != io_in_bits_1_bp_br_taken | _bp_wrong_T_13; // @[EXU.scala 131:58]
  wire  _bp_wrong_T_15 = _bp_wrong_T_14 & io_in_valid; // @[EXU.scala 132:131]
  wire  _bp_wrong_T_5 = br_taken & io_in_bits_0_bp_br_taken & (br_target != io_in_bits_0_bp_br_target | br_type !=
    io_in_bits_0_bp_br_type); // @[EXU.scala 132:45]
  wire  _bp_wrong_T_6 = br_taken != io_in_bits_0_bp_br_taken | _bp_wrong_T_5; // @[EXU.scala 131:58]
  wire  _bp_wrong_T_7 = _bp_wrong_T_6 & io_in_valid; // @[EXU.scala 132:131]
  wire  _GEN_37 = _T_5 & _bp_wrong_T_7; // @[EXU.scala 121:62 EXU.scala 131:16 EXU.scala 119:12]
  wire  bp_wrong = _T_7 ? _bp_wrong_T_15 : _GEN_37; // @[EXU.scala 121:62 EXU.scala 131:16]
  wire  _frontend_reflush_T_4 = (csr_is_reflush & ~handle_int | fence | bp_wrong) & io_in_valid; // @[EXU.scala 228:79]
  reg  frontend_reflush_reg; // @[EXU.scala 222:37]
  wire  _frontend_reflush_T_6 = frontend_reflush_reg & io_out_valid; // @[EXU.scala 229:26]
  wire  _frontend_reflush_T_7 = (csr_is_reflush & ~handle_int | fence | bp_wrong) & io_in_valid & io_out_valid |
    _frontend_reflush_T_6; // @[EXU.scala 228:111]
  wire  frontend_reflush = _frontend_reflush_T_7 | handle_int; // @[EXU.scala 229:42]
  wire  _GEN_28 = _T_5 & io_in_valid; // @[EXU.scala 121:62 EXU.scala 122:20 EXU.scala 117:10]
  wire  _GEN_30 = _T_5 & br_taken; // @[EXU.scala 121:62 EXU.scala 124:23 EXU.scala 117:10]
  wire [31:0] _GEN_31 = _T_5 ? br_target : 32'h0; // @[EXU.scala 121:62 EXU.scala 125:24 EXU.scala 117:10]
  wire [1:0] _GEN_32 = _T_5 ? br_type : 2'h0; // @[EXU.scala 121:62 EXU.scala 126:22 EXU.scala 117:10]
  wire  _GEN_33 = _T_5 & bp_wrong; // @[EXU.scala 121:62 EXU.scala 127:23 EXU.scala 117:10]
  wire [2:0] _GEN_35 = _T_5 ? call_count : 3'h0; // @[EXU.scala 121:62 EXU.scala 129:25 EXU.scala 117:10]
  wire [2:0] _GEN_36 = _T_5 ? ret_count : 3'h0; // @[EXU.scala 121:62 EXU.scala 130:24 EXU.scala 117:10]
  wire  is_clint = (clint_io_is_mtime | clint_io_is_mtimecmp) & io_in_valid; // @[EXU.scala 192:59]
  wire [63:0] lsu_rdata = is_clint ? clint_io_rdata : lsu_io_rdata; // @[EXU.scala 149:19]
  wire  _T_17 = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid; // @[EXU.scala 151:41]
  wire  _GEN_48 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid & io_in_valid; // @[EXU.scala 151:62 EXU.scala 152:14 EXU.scala 138:10]
  wire  is_lsu = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? io_in_valid : _GEN_48; // @[EXU.scala 151:62 EXU.scala 152:14]
  wire  _lsu_io_is_lsu_T_1 = is_lsu & ~is_clint; // @[EXU.scala 156:31]
  wire [63:0] _GEN_49 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid ? io_in_bits_0_src1_value : 64'h0; // @[EXU.scala 151:62 EXU.scala 153:19 EXU.scala 139:15]
  wire [63:0] _GEN_50 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid ? io_in_bits_0_src2_value : 64'h0; // @[EXU.scala 151:62 EXU.scala 154:19 EXU.scala 140:15]
  wire [63:0] _GEN_51 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid ? io_in_bits_0_rs2_value : 64'h0; // @[EXU.scala 151:62 EXU.scala 155:20 EXU.scala 141:16]
  wire  _GEN_52 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid & (is_lsu & ~is_clint); // @[EXU.scala 151:62 EXU.scala 156:21 EXU.scala 142:17]
  wire  _GEN_53 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid & io_in_bits_0_wen; // @[EXU.scala 151:62 EXU.scala 157:18 EXU.scala 143:14]
  wire [3:0] _GEN_54 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid ? io_in_bits_0_lsu_op : 4'h0; // @[EXU.scala 151:62 EXU.scala 158:21 EXU.scala 144:17]
  wire  _GEN_55 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid & is_mdu; // @[EXU.scala 151:62 EXU.scala 159:21 EXU.scala 145:17]
  wire  mdu_ok = mdu_io_result_ok;
  wire  _GEN_56 = io_in_bits_0_fu_type == 3'h2 & io_in_bits_0_valid & mdu_ok; // @[EXU.scala 151:62 EXU.scala 160:21 EXU.scala 146:17]
  wire [2:0] _csr_io_csr_op_T_1 = io_in_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [2:0] _csr_io_csr_op_T_2 = io_in_bits_0_csr_op & _csr_io_csr_op_T_1; // @[EXU.scala 179:42]
  wire [31:0] _GEN_66 = io_in_bits_0_fu_type == 3'h3 & io_in_bits_0_valid ? io_in_bits_0_pc : 32'h0; // @[EXU.scala 177:62 EXU.scala 178:17 EXU.scala 165:13]
  wire [2:0] _GEN_67 = io_in_bits_0_fu_type == 3'h3 & io_in_bits_0_valid ? _csr_io_csr_op_T_2 : 3'h0; // @[EXU.scala 177:62 EXU.scala 179:21 EXU.scala 166:17]
  wire [11:0] _GEN_68 = io_in_bits_0_fu_type == 3'h3 & io_in_bits_0_valid ? io_in_bits_0_inst[31:20] : 12'h0; // @[EXU.scala 177:62 EXU.scala 180:19 EXU.scala 167:15]
  wire [63:0] _GEN_69 = io_in_bits_0_fu_type == 3'h3 & io_in_bits_0_valid ? io_in_bits_0_src1_value : 64'h0; // @[EXU.scala 177:62 EXU.scala 181:18 EXU.scala 168:14]
  wire  _GEN_70 = io_in_bits_0_fu_type == 3'h3 & io_in_bits_0_valid & io_in_valid; // @[EXU.scala 177:62 EXU.scala 182:20 EXU.scala 169:16]
  wire [2:0] _csr_io_csr_op_T_5 = io_in_bits_1_csr_op & _csr_io_csr_op_T_1; // @[EXU.scala 179:42]
  wire [31:0] lsu_addr = lsu_io_addr; // @[EXU.scala 34:22 EXU.scala 148:12]
  wire [63:0] _GEN_108 = {{32'd0}, lsu_addr}; // @[EXU.scala 189:34]
  wire [31:0] _final_result_0_T_1 = io_in_bits_0_pc + 32'h4; // @[EXU.scala 204:32]
  wire [63:0] alu_result_0 = alu_0_io_result;
  wire [63:0] _final_result_0_T_3 = 3'h0 == io_in_bits_0_fu_type ? alu_result_0 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] mdu_result = mdu_io_result;
  wire [63:0] _final_result_0_T_5 = 3'h4 == io_in_bits_0_fu_type ? mdu_result : _final_result_0_T_3; // @[Mux.scala 80:57]
  wire [63:0] _final_result_0_T_7 = 3'h1 == io_in_bits_0_fu_type ? {{32'd0}, _final_result_0_T_1} : _final_result_0_T_5; // @[Mux.scala 80:57]
  wire [63:0] _final_result_0_T_9 = 3'h2 == io_in_bits_0_fu_type ? lsu_rdata : _final_result_0_T_7; // @[Mux.scala 80:57]
  wire [63:0] csr_rdata = csr_io_rdata; // @[EXU.scala 36:23 EXU.scala 170:13]
  wire [31:0] _final_result_1_T_1 = io_in_bits_1_pc + 32'h4; // @[EXU.scala 204:32]
  wire [63:0] alu_result_1 = alu_1_io_result;
  wire [63:0] _final_result_1_T_3 = 3'h0 == io_in_bits_1_fu_type ? alu_result_1 : 64'h0; // @[Mux.scala 80:57]
  wire [63:0] _final_result_1_T_5 = 3'h4 == io_in_bits_1_fu_type ? mdu_result : _final_result_1_T_3; // @[Mux.scala 80:57]
  wire [63:0] _final_result_1_T_7 = 3'h1 == io_in_bits_1_fu_type ? {{32'd0}, _final_result_1_T_1} : _final_result_1_T_5; // @[Mux.scala 80:57]
  wire [63:0] _final_result_1_T_9 = 3'h2 == io_in_bits_1_fu_type ? lsu_rdata : _final_result_1_T_7; // @[Mux.scala 80:57]
  wire  _T_33 = 2'h0 == blk_state; // @[Conditional.scala 37:30]
  wire  _GEN_82 = is_mdu ? 1'h0 : 1'h1; // @[EXU.scala 240:28 EXU.scala 241:19 EXU.scala 233:17]
  wire  _GEN_84 = _lsu_io_is_lsu_T_1 ? 1'h0 : _GEN_82; // @[EXU.scala 237:41 EXU.scala 238:19]
  wire  _GEN_86 = _lsu_io_is_lsu_T_1 & is_mdu ? 1'h0 : _GEN_84; // @[EXU.scala 234:46 EXU.scala 235:19]
  wire  _T_39 = 2'h3 == blk_state; // @[Conditional.scala 37:30]
  wire  _T_40 = io_dmem_data_ok & mdu_ok; // @[EXU.scala 247:29]
  wire  _T_41 = 2'h1 == blk_state; // @[Conditional.scala 37:30]
  wire  _T_42 = 2'h2 == blk_state; // @[Conditional.scala 37:30]
  wire  _GEN_96 = _T_42 ? io_dmem_data_ok : 1'h1; // @[Conditional.scala 39:67]
  wire  _GEN_98 = _T_41 ? mdu_ok : _GEN_96; // @[Conditional.scala 39:67]
  wire  _GEN_100 = _T_39 ? _T_40 : _GEN_98; // @[Conditional.scala 39:67]
  wire  blk_ready = _T_33 ? _GEN_86 : _GEN_100; // @[Conditional.scala 40:58]
  wire  _GEN_80 = io_out_valid ? 1'h0 : frontend_reflush_reg; // @[EXU.scala 225:30 EXU.scala 226:26 EXU.scala 222:37]
  wire  _GEN_81 = _frontend_reflush_T_4 & ~io_out_valid | _GEN_80; // @[EXU.scala 223:97 EXU.scala 224:26]
  wire [1:0] _GEN_83 = is_mdu ? 2'h1 : blk_state; // @[EXU.scala 240:28 EXU.scala 242:19 EXU.scala 51:26]
  wire [1:0] _GEN_88 = mdu_ok ? 2'h2 : blk_state; // @[EXU.scala 252:28 EXU.scala 253:19 EXU.scala 51:26]
  wire [1:0] _GEN_89 = io_dmem_data_ok ? 2'h1 : _GEN_88; // @[EXU.scala 250:37 EXU.scala 251:19]
  wire [1:0] _GEN_93 = mdu_ok ? 2'h0 : blk_state; // @[EXU.scala 258:21 EXU.scala 260:19 EXU.scala 51:26]
  wire [1:0] _GEN_95 = io_dmem_data_ok ? 2'h0 : blk_state; // @[EXU.scala 265:29 EXU.scala 267:19 EXU.scala 51:26]
  wire [1:0] _GEN_97 = _T_42 ? _GEN_95 : blk_state; // @[Conditional.scala 39:67 EXU.scala 51:26]
  wire [31:0] _GEN_104 = (_T_4 | fence) & io_in_bits_0_valid ? _final_result_0_T_1 : 32'h0; // @[EXU.scala 281:73 EXU.scala 282:22]
  wire [31:0] static_next_pc = (_T_6 | fence) & io_in_bits_1_valid ? _final_result_1_T_1 : _GEN_104; // @[EXU.scala 281:73 EXU.scala 282:22]
  wire [31:0] _io_reflush_bus_br_target_T_1 = bp_wrong & br_taken ? br_target : static_next_pc; // @[EXU.scala 287:8]
  wire [31:0] csr_target = csr_io_csr_target; // @[EXU.scala 44:24 EXU.scala 172:14]
  ALU alu_0 ( // @[EXU.scala 20:21]
    .io_alu_op(alu_0_io_alu_op),
    .io_rv64(alu_0_io_rv64),
    .io_src1(alu_0_io_src1),
    .io_src2(alu_0_io_src2),
    .io_result(alu_0_io_result)
  );
  ALU alu_1 ( // @[EXU.scala 20:21]
    .io_alu_op(alu_1_io_alu_op),
    .io_rv64(alu_1_io_rv64),
    .io_src1(alu_1_io_src1),
    .io_src2(alu_1_io_src2),
    .io_result(alu_1_io_result)
  );
  MDU mdu ( // @[EXU.scala 23:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_mdu_op(mdu_io_mdu_op),
    .io_rv64(mdu_io_rv64),
    .io_src1(mdu_io_src1),
    .io_src2(mdu_io_src2),
    .io_result_ok(mdu_io_result_ok),
    .io_result(mdu_io_result)
  );
  BRU bru ( // @[EXU.scala 24:19]
    .io_bru_op(bru_io_bru_op),
    .io_src1(bru_io_src1),
    .io_src2(bru_io_src2),
    .io_pc(bru_io_pc),
    .io_imm(bru_io_imm),
    .io_br_taken(bru_io_br_taken),
    .io_br_target(bru_io_br_target),
    .io_rs1(bru_io_rs1),
    .io_rd(bru_io_rd),
    .io_btb_type(bru_io_btb_type)
  );
  LSU lsu ( // @[EXU.scala 25:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_dmem_valid(lsu_io_dmem_valid),
    .io_dmem_op(lsu_io_dmem_op),
    .io_dmem_addr(lsu_io_dmem_addr),
    .io_dmem_wstrb(lsu_io_dmem_wstrb),
    .io_dmem_wdata(lsu_io_dmem_wdata),
    .io_dmem_fence(lsu_io_dmem_fence),
    .io_dmem_fence_finish(lsu_io_dmem_fence_finish),
    .io_dmem_data_ok(lsu_io_dmem_data_ok),
    .io_dmem_rdata(lsu_io_dmem_rdata),
    .io_src1(lsu_io_src1),
    .io_src2(lsu_io_src2),
    .io_wdata(lsu_io_wdata),
    .io_addr(lsu_io_addr),
    .io_is_lsu(lsu_io_is_lsu),
    .io_wen(lsu_io_wen),
    .io_lsu_op(lsu_io_lsu_op),
    .io_rdata(lsu_io_rdata),
    .io_is_mdu(lsu_io_is_mdu),
    .io_mdu_ok(lsu_io_mdu_ok),
    .dcache_fence_finish_0(lsu_dcache_fence_finish_0),
    .fence_i(lsu_fence_i),
    .icache_fence_finish_0(lsu_icache_fence_finish_0)
  );
  CSR csr ( // @[EXU.scala 26:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_pc(csr_io_pc),
    .io_csr_op(csr_io_csr_op),
    .io_addr(csr_io_addr),
    .io_src(csr_io_src),
    .io_rdata(csr_io_rdata),
    .io_is_reflush(csr_io_is_reflush),
    .io_csr_target(csr_io_csr_target),
    .io_handle_int(csr_io_handle_int),
    .io_valid(csr_io_valid),
    .clint_has_int(csr_clint_has_int)
  );
  CLINT clint ( // @[EXU.scala 27:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io_is_mtime(clint_io_is_mtime),
    .io_is_mtimecmp(clint_io_is_mtimecmp),
    .io_is_clint(clint_io_is_clint),
    .io_wen(clint_io_wen),
    .io_wdata(clint_io_wdata),
    .io_rdata(clint_io_rdata),
    .has_int_0(clint_has_int_0)
  );
  assign io_dmem_valid = lsu_io_dmem_valid; // @[EXU.scala 147:15]
  assign io_dmem_op = lsu_io_dmem_op; // @[EXU.scala 147:15]
  assign io_dmem_addr = lsu_io_dmem_addr; // @[EXU.scala 147:15]
  assign io_dmem_wstrb = lsu_io_dmem_wstrb; // @[EXU.scala 147:15]
  assign io_dmem_wdata = lsu_io_dmem_wdata; // @[EXU.scala 147:15]
  assign io_dmem_fence = lsu_io_dmem_fence; // @[EXU.scala 147:15]
  assign io_in_ready = blk_ready | ~io_in_valid; // @[EXU.scala 220:46]
  assign io_out_valid = io_in_valid & _frontend_reflush_T & blk_ready; // @[EXU.scala 219:46]
  assign io_out_bits_0_valid = io_in_bits_0_valid; // @[EXU.scala 211:26]
  assign io_out_bits_0_pc = io_in_bits_0_pc; // @[EXU.scala 212:23]
  assign io_out_bits_0_final_result = 3'h3 == io_in_bits_0_fu_type ? csr_rdata : _final_result_0_T_9; // @[Mux.scala 80:57]
  assign io_out_bits_0_dest = io_in_bits_0_dest; // @[EXU.scala 215:25]
  assign io_out_bits_0_wen = io_in_bits_0_wen; // @[EXU.scala 216:24]
  assign io_out_bits_1_valid = io_in_bits_1_valid; // @[EXU.scala 211:26]
  assign io_out_bits_1_final_result = 3'h3 == io_in_bits_1_fu_type ? csr_rdata : _final_result_1_T_9; // @[Mux.scala 80:57]
  assign io_out_bits_1_dest = io_in_bits_1_dest; // @[EXU.scala 215:25]
  assign io_out_bits_1_wen = io_in_bits_1_wen; // @[EXU.scala 216:24]
  assign io_forward_0_blk_valid = io_forward_0_fwd_valid & ~blk_ready; // @[EXU.scala 272:56]
  assign io_forward_0_fwd_valid = io_in_bits_0_wen & io_in_bits_0_dest != 5'h0 & io_in_valid & io_in_bits_0_valid; // @[EXU.scala 273:89]
  assign io_forward_0_rf_waddr = io_in_bits_0_dest; // @[EXU.scala 274:28]
  assign io_forward_0_rf_wdata = 3'h3 == io_in_bits_0_fu_type ? csr_rdata : _final_result_0_T_9; // @[Mux.scala 80:57]
  assign io_forward_1_blk_valid = io_forward_1_fwd_valid & ~blk_ready; // @[EXU.scala 272:56]
  assign io_forward_1_fwd_valid = io_in_bits_1_wen & io_in_bits_1_dest != 5'h0 & io_in_valid & io_in_bits_1_valid; // @[EXU.scala 273:89]
  assign io_forward_1_rf_waddr = io_in_bits_1_dest; // @[EXU.scala 274:28]
  assign io_forward_1_rf_wdata = 3'h3 == io_in_bits_1_fu_type ? csr_rdata : _final_result_1_T_9; // @[Mux.scala 80:57]
  assign io_reflush_bus_is_reflush = frontend_reflush; // @[EXU.scala 278:29]
  assign io_reflush_bus_br_target = csr_is_reflush ? csr_target : _io_reflush_bus_br_target_T_1; // @[EXU.scala 286:34]
  assign io_bpu_valid = _T_7 ? io_in_valid : _GEN_28; // @[EXU.scala 121:62 EXU.scala 122:20]
  assign io_bpu_pc = _T_7 ? io_in_bits_1_pc : _GEN_13; // @[EXU.scala 121:62 EXU.scala 123:17]
  assign io_bpu_bp_taken = _T_7 ? br_taken : _GEN_30; // @[EXU.scala 121:62 EXU.scala 124:23]
  assign io_bpu_bp_target = _T_7 ? br_target : _GEN_31; // @[EXU.scala 121:62 EXU.scala 125:24]
  assign io_bpu_bp_type = _T_7 ? br_type : _GEN_32; // @[EXU.scala 121:62 EXU.scala 126:22]
  assign io_bpu_bp_wrong = _T_7 ? bp_wrong : _GEN_33; // @[EXU.scala 121:62 EXU.scala 127:23]
  assign io_bpu_fence = fence; // @[EXU.scala 118:16]
  assign io_bpu_call_count = _T_7 ? call_count : _GEN_35; // @[EXU.scala 121:62 EXU.scala 129:25]
  assign io_bpu_ret_count = _T_7 ? ret_count : _GEN_36; // @[EXU.scala 121:62 EXU.scala 130:24]
  assign frontend_reflush_0 = frontend_reflush;
  assign dcache_fence_finish = lsu_dcache_fence_finish_0;
  assign fence_0 = fence;
  assign alu_0_io_alu_op = io_in_bits_0_alu_op; // @[EXU.scala 57:22]
  assign alu_0_io_rv64 = io_in_bits_0_rv64; // @[EXU.scala 58:20]
  assign alu_0_io_src1 = io_in_bits_0_src1_value; // @[EXU.scala 59:20]
  assign alu_0_io_src2 = io_in_bits_0_src2_value; // @[EXU.scala 60:20]
  assign alu_1_io_alu_op = io_in_bits_1_alu_op; // @[EXU.scala 57:22]
  assign alu_1_io_rv64 = io_in_bits_1_rv64; // @[EXU.scala 58:20]
  assign alu_1_io_src1 = io_in_bits_1_src1_value; // @[EXU.scala 59:20]
  assign alu_1_io_src2 = io_in_bits_1_src2_value; // @[EXU.scala 60:20]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_mdu_op = io_in_bits_1_fu_type == 3'h4 & io_in_bits_1_valid ? _mdu_io_mdu_op_T_5 : _GEN_3; // @[EXU.scala 72:61 EXU.scala 76:21]
  assign mdu_io_rv64 = io_in_bits_1_fu_type == 3'h4 & io_in_bits_1_valid ? io_in_bits_1_rv64 : _GEN_4; // @[EXU.scala 72:61 EXU.scala 77:19]
  assign mdu_io_src1 = io_in_bits_1_fu_type == 3'h4 & io_in_bits_1_valid ? io_in_bits_1_src1_value : _GEN_1; // @[EXU.scala 72:61 EXU.scala 74:19]
  assign mdu_io_src2 = io_in_bits_1_fu_type == 3'h4 & io_in_bits_1_valid ? io_in_bits_1_src2_value : _GEN_2; // @[EXU.scala 72:61 EXU.scala 75:19]
  assign bru_io_bru_op = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_bru_op : _GEN_10; // @[EXU.scala 94:62 EXU.scala 95:21]
  assign bru_io_src1 = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_src1_value : _GEN_11; // @[EXU.scala 94:62 EXU.scala 96:19]
  assign bru_io_src2 = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_src2_value : _GEN_12; // @[EXU.scala 94:62 EXU.scala 97:19]
  assign bru_io_pc = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_pc : _GEN_13; // @[EXU.scala 94:62 EXU.scala 98:17]
  assign bru_io_imm = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_imm : _GEN_14; // @[EXU.scala 94:62 EXU.scala 99:18]
  assign bru_io_rs1 = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_rs1 : _GEN_15; // @[EXU.scala 94:62 EXU.scala 100:18]
  assign bru_io_rd = io_in_bits_1_fu_type == 3'h1 & io_in_bits_1_valid ? io_in_bits_1_dest : _GEN_16; // @[EXU.scala 94:62 EXU.scala 101:17]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_dmem_fence_finish = io_dmem_fence_finish; // @[EXU.scala 147:15]
  assign lsu_io_dmem_data_ok = io_dmem_data_ok; // @[EXU.scala 147:15]
  assign lsu_io_dmem_rdata = io_dmem_rdata; // @[EXU.scala 147:15]
  assign lsu_io_src1 = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? io_in_bits_1_src1_value : _GEN_49; // @[EXU.scala 151:62 EXU.scala 153:19]
  assign lsu_io_src2 = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? io_in_bits_1_src2_value : _GEN_50; // @[EXU.scala 151:62 EXU.scala 154:19]
  assign lsu_io_wdata = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? io_in_bits_1_rs2_value : _GEN_51; // @[EXU.scala 151:62 EXU.scala 155:20]
  assign lsu_io_is_lsu = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? is_lsu & ~is_clint : _GEN_52; // @[EXU.scala 151:62 EXU.scala 156:21]
  assign lsu_io_wen = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? io_in_bits_1_wen : _GEN_53; // @[EXU.scala 151:62 EXU.scala 157:18]
  assign lsu_io_lsu_op = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? io_in_bits_1_lsu_op : _GEN_54; // @[EXU.scala 151:62 EXU.scala 158:21]
  assign lsu_io_is_mdu = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? is_mdu : _GEN_55; // @[EXU.scala 151:62 EXU.scala 159:21]
  assign lsu_io_mdu_ok = io_in_bits_1_fu_type == 3'h2 & io_in_bits_1_valid ? mdu_ok : _GEN_56; // @[EXU.scala 151:62 EXU.scala 160:21]
  assign lsu_fence_i = fence_0;
  assign lsu_icache_fence_finish_0 = icache_fence_finish;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_pc = io_in_bits_1_fu_type == 3'h3 & io_in_bits_1_valid ? io_in_bits_1_pc : _GEN_66; // @[EXU.scala 177:62 EXU.scala 178:17]
  assign csr_io_csr_op = io_in_bits_1_fu_type == 3'h3 & io_in_bits_1_valid ? _csr_io_csr_op_T_5 : _GEN_67; // @[EXU.scala 177:62 EXU.scala 179:21]
  assign csr_io_addr = io_in_bits_1_fu_type == 3'h3 & io_in_bits_1_valid ? io_in_bits_1_inst[31:20] : _GEN_68; // @[EXU.scala 177:62 EXU.scala 180:19]
  assign csr_io_src = io_in_bits_1_fu_type == 3'h3 & io_in_bits_1_valid ? io_in_bits_1_src1_value : _GEN_69; // @[EXU.scala 177:62 EXU.scala 181:18]
  assign csr_io_valid = io_in_bits_1_fu_type == 3'h3 & io_in_bits_1_valid ? io_in_valid : _GEN_70; // @[EXU.scala 177:62 EXU.scala 182:20]
  assign csr_clint_has_int = clint_has_int_0;
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io_is_mtime = _GEN_108 == 64'h200bff8; // @[EXU.scala 189:34]
  assign clint_io_is_mtimecmp = _GEN_108 == 64'h2004000; // @[EXU.scala 190:37]
  assign clint_io_is_clint = is_lsu & is_clint; // @[EXU.scala 191:31]
  assign clint_io_wen = _T_17 ? io_in_bits_1_wen : _GEN_53; // @[EXU.scala 194:62 EXU.scala 195:20]
  assign clint_io_wdata = _T_17 ? io_in_bits_1_rs2_value : _GEN_51; // @[EXU.scala 194:62 EXU.scala 196:22]
  always @(posedge clock) begin
    if (reset) begin // @[EXU.scala 51:26]
      blk_state <= 2'h0; // @[EXU.scala 51:26]
    end else if (_T_33) begin // @[Conditional.scala 40:58]
      if (_lsu_io_is_lsu_T_1 & is_mdu) begin // @[EXU.scala 234:46]
        blk_state <= 2'h3; // @[EXU.scala 236:19]
      end else if (_lsu_io_is_lsu_T_1) begin // @[EXU.scala 237:41]
        blk_state <= 2'h2; // @[EXU.scala 239:19]
      end else begin
        blk_state <= _GEN_83;
      end
    end else if (_T_39) begin // @[Conditional.scala 39:67]
      if (io_dmem_data_ok & mdu_ok) begin // @[EXU.scala 247:40]
        blk_state <= 2'h0; // @[EXU.scala 249:19]
      end else begin
        blk_state <= _GEN_89;
      end
    end else if (_T_41) begin // @[Conditional.scala 39:67]
      blk_state <= _GEN_93;
    end else begin
      blk_state <= _GEN_97;
    end
    if (reset) begin // @[EXU.scala 106:27]
      call_count <= 3'h0; // @[EXU.scala 106:27]
    end else if (frontend_reflush) begin // @[EXU.scala 109:27]
      call_count <= 3'h0; // @[EXU.scala 110:16]
    end else if (io_bpu_valid & blk_state == 2'h0) begin // @[EXU.scala 112:56]
      call_count <= _call_count_T_2; // @[EXU.scala 113:16]
    end
    if (reset) begin // @[EXU.scala 107:26]
      ret_count <= 3'h0; // @[EXU.scala 107:26]
    end else if (frontend_reflush) begin // @[EXU.scala 109:27]
      ret_count <= 3'h0; // @[EXU.scala 111:15]
    end else if (io_bpu_valid & blk_state == 2'h0) begin // @[EXU.scala 112:56]
      ret_count <= _ret_count_T_2; // @[EXU.scala 114:15]
    end
    if (reset) begin // @[EXU.scala 222:37]
      frontend_reflush_reg <= 1'h0; // @[EXU.scala 222:37]
    end else begin
      frontend_reflush_reg <= _GEN_81;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  blk_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  call_count = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  ret_count = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  frontend_reflush_reg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         io__in_valid,
  input         io__in_bits_0_valid,
  input  [31:0] io__in_bits_0_pc,
  input  [63:0] io__in_bits_0_final_result,
  input  [4:0]  io__in_bits_0_dest,
  input         io__in_bits_0_wen,
  input         io__in_bits_1_valid,
  input  [63:0] io__in_bits_1_final_result,
  input  [4:0]  io__in_bits_1_dest,
  input         io__in_bits_1_wen,
  output        io__wb_bus_0_rf_wen,
  output [4:0]  io__wb_bus_0_rf_waddr,
  output [63:0] io__wb_bus_0_rf_wdata,
  output        io__wb_bus_1_rf_wen,
  output [4:0]  io__wb_bus_1_rf_waddr,
  output [63:0] io__wb_bus_1_rf_wdata,
  output [31:0] io__commit_0_pc,
  output [31:0] io_commit_0_pc
);
  assign io__wb_bus_0_rf_wen = io__in_bits_0_wen & io__in_bits_0_dest != 5'h0 & io__in_valid & io__in_bits_0_valid; // @[WBU.scala 17:85]
  assign io__wb_bus_0_rf_waddr = io__in_bits_0_dest; // @[WBU.scala 18:27]
  assign io__wb_bus_0_rf_wdata = io__in_bits_0_final_result; // @[WBU.scala 19:27]
  assign io__wb_bus_1_rf_wen = io__in_bits_1_wen & io__in_bits_1_dest != 5'h0 & io__in_valid & io__in_bits_1_valid; // @[WBU.scala 17:85]
  assign io__wb_bus_1_rf_waddr = io__in_bits_1_dest; // @[WBU.scala 18:27]
  assign io__wb_bus_1_rf_wdata = io__in_bits_1_final_result; // @[WBU.scala 19:27]
  assign io__commit_0_pc = io__in_bits_0_pc; // @[WBU.scala 21:21]
  assign io_commit_0_pc = io__commit_0_pc;
endmodule
module BTB(
  input         clock,
  input         reset,
  input         io_wen,
  input  [2:0]  io_index_r,
  input  [2:0]  io_index_w,
  input  [24:0] io_in_tag,
  input  [1:0]  io_in_offset,
  input  [1:0]  io_in_btb_type,
  input  [31:0] io_in_target,
  output [24:0] io_out_tag,
  output [1:0]  io_out_offset,
  output [1:0]  io_out_btb_type,
  output [31:0] io_out_target,
  output        io_valid_r,
  input         io_fence
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
`endif // RANDOMIZE_REG_INIT
  reg [24:0] btb_entry_0_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_0_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_0_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_0_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_1_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_1_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_1_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_1_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_2_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_2_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_2_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_2_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_3_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_3_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_3_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_3_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_4_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_4_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_4_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_4_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_5_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_5_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_5_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_5_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_6_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_6_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_6_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_6_target; // @[BPU.scala 33:26]
  reg [24:0] btb_entry_7_tag; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_7_offset; // @[BPU.scala 33:26]
  reg [1:0] btb_entry_7_btb_type; // @[BPU.scala 33:26]
  reg [31:0] btb_entry_7_target; // @[BPU.scala 33:26]
  reg  valid_0; // @[BPU.scala 34:22]
  reg  valid_1; // @[BPU.scala 34:22]
  reg  valid_2; // @[BPU.scala 34:22]
  reg  valid_3; // @[BPU.scala 34:22]
  reg  valid_4; // @[BPU.scala 34:22]
  reg  valid_5; // @[BPU.scala 34:22]
  reg  valid_6; // @[BPU.scala 34:22]
  reg  valid_7; // @[BPU.scala 34:22]
  wire  _GEN_32 = 3'h0 == io_index_w | valid_0; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_33 = 3'h1 == io_index_w | valid_1; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_34 = 3'h2 == io_index_w | valid_2; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_35 = 3'h3 == io_index_w | valid_3; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_36 = 3'h4 == io_index_w | valid_4; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_37 = 3'h5 == io_index_w | valid_5; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_38 = 3'h6 == io_index_w | valid_6; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  wire  _GEN_39 = 3'h7 == io_index_w | valid_7; // @[BPU.scala 41:20 BPU.scala 41:20 BPU.scala 34:22]
  reg [24:0] io_out_tag_REG; // @[BPU.scala 44:21]
  wire [24:0] _GEN_81 = 3'h1 == io_index_r ? btb_entry_1_tag : btb_entry_0_tag; // @[BPU.scala 44:21 BPU.scala 44:21]
  wire [24:0] _GEN_82 = 3'h2 == io_index_r ? btb_entry_2_tag : _GEN_81; // @[BPU.scala 44:21 BPU.scala 44:21]
  wire [24:0] _GEN_83 = 3'h3 == io_index_r ? btb_entry_3_tag : _GEN_82; // @[BPU.scala 44:21 BPU.scala 44:21]
  wire [24:0] _GEN_84 = 3'h4 == io_index_r ? btb_entry_4_tag : _GEN_83; // @[BPU.scala 44:21 BPU.scala 44:21]
  reg [1:0] io_out_offset_REG; // @[BPU.scala 45:24]
  wire [1:0] _GEN_89 = 3'h1 == io_index_r ? btb_entry_1_offset : btb_entry_0_offset; // @[BPU.scala 45:24 BPU.scala 45:24]
  wire [1:0] _GEN_90 = 3'h2 == io_index_r ? btb_entry_2_offset : _GEN_89; // @[BPU.scala 45:24 BPU.scala 45:24]
  wire [1:0] _GEN_91 = 3'h3 == io_index_r ? btb_entry_3_offset : _GEN_90; // @[BPU.scala 45:24 BPU.scala 45:24]
  wire [1:0] _GEN_92 = 3'h4 == io_index_r ? btb_entry_4_offset : _GEN_91; // @[BPU.scala 45:24 BPU.scala 45:24]
  reg [31:0] io_out_target_REG; // @[BPU.scala 46:24]
  wire [31:0] _GEN_97 = 3'h1 == io_index_r ? btb_entry_1_target : btb_entry_0_target; // @[BPU.scala 46:24 BPU.scala 46:24]
  wire [31:0] _GEN_98 = 3'h2 == io_index_r ? btb_entry_2_target : _GEN_97; // @[BPU.scala 46:24 BPU.scala 46:24]
  wire [31:0] _GEN_99 = 3'h3 == io_index_r ? btb_entry_3_target : _GEN_98; // @[BPU.scala 46:24 BPU.scala 46:24]
  wire [31:0] _GEN_100 = 3'h4 == io_index_r ? btb_entry_4_target : _GEN_99; // @[BPU.scala 46:24 BPU.scala 46:24]
  reg [1:0] io_out_btb_type_REG; // @[BPU.scala 47:26]
  wire [1:0] _GEN_105 = 3'h1 == io_index_r ? btb_entry_1_btb_type : btb_entry_0_btb_type; // @[BPU.scala 47:26 BPU.scala 47:26]
  wire [1:0] _GEN_106 = 3'h2 == io_index_r ? btb_entry_2_btb_type : _GEN_105; // @[BPU.scala 47:26 BPU.scala 47:26]
  wire [1:0] _GEN_107 = 3'h3 == io_index_r ? btb_entry_3_btb_type : _GEN_106; // @[BPU.scala 47:26 BPU.scala 47:26]
  wire [1:0] _GEN_108 = 3'h4 == io_index_r ? btb_entry_4_btb_type : _GEN_107; // @[BPU.scala 47:26 BPU.scala 47:26]
  reg  io_valid_r_REG; // @[BPU.scala 48:24]
  wire  _GEN_113 = 3'h1 == io_index_r ? valid_1 : valid_0; // @[BPU.scala 48:24 BPU.scala 48:24]
  wire  _GEN_114 = 3'h2 == io_index_r ? valid_2 : _GEN_113; // @[BPU.scala 48:24 BPU.scala 48:24]
  wire  _GEN_115 = 3'h3 == io_index_r ? valid_3 : _GEN_114; // @[BPU.scala 48:24 BPU.scala 48:24]
  wire  _GEN_116 = 3'h4 == io_index_r ? valid_4 : _GEN_115; // @[BPU.scala 48:24 BPU.scala 48:24]
  assign io_out_tag = io_out_tag_REG; // @[BPU.scala 44:11]
  assign io_out_offset = io_out_offset_REG; // @[BPU.scala 45:14]
  assign io_out_btb_type = io_out_btb_type_REG; // @[BPU.scala 47:16]
  assign io_out_target = io_out_target_REG; // @[BPU.scala 46:14]
  assign io_valid_r = io_valid_r_REG; // @[BPU.scala 48:14]
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_0_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h0 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_0_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_0_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h0 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_0_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_0_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h0 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_0_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_0_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h0 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_0_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_1_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h1 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_1_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_1_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h1 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_1_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_1_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h1 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_1_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_1_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h1 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_1_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_2_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h2 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_2_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_2_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h2 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_2_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_2_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h2 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_2_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_2_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h2 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_2_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_3_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h3 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_3_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_3_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h3 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_3_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_3_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h3 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_3_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_3_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h3 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_3_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_4_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h4 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_4_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_4_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h4 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_4_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_4_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h4 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_4_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_4_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h4 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_4_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_5_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h5 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_5_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_5_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h5 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_5_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_5_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h5 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_5_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_5_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h5 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_5_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_6_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h6 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_6_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_6_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h6 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_6_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_6_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h6 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_6_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_6_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h6 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_6_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_7_tag <= 25'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h7 == io_index_w) begin // @[BPU.scala 37:28]
        btb_entry_7_tag <= io_in_tag; // @[BPU.scala 37:28]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_7_offset <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h7 == io_index_w) begin // @[BPU.scala 38:31]
        btb_entry_7_offset <= io_in_offset; // @[BPU.scala 38:31]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_7_btb_type <= 2'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h7 == io_index_w) begin // @[BPU.scala 40:33]
        btb_entry_7_btb_type <= io_in_btb_type; // @[BPU.scala 40:33]
      end
    end
    if (reset) begin // @[BPU.scala 33:26]
      btb_entry_7_target <= 32'h0; // @[BPU.scala 33:26]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      if (3'h7 == io_index_w) begin // @[BPU.scala 39:31]
        btb_entry_7_target <= io_in_target; // @[BPU.scala 39:31]
      end
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_0 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_0 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_0 <= _GEN_32;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_1 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_1 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_1 <= _GEN_33;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_2 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_2 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_2 <= _GEN_34;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_3 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_3 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_3 <= _GEN_35;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_4 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_4 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_4 <= _GEN_36;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_5 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_5 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_5 <= _GEN_37;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_6 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_6 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_6 <= _GEN_38;
    end
    if (reset) begin // @[BPU.scala 34:22]
      valid_7 <= 1'h0; // @[BPU.scala 34:22]
    end else if (reset | io_fence) begin // @[BPU.scala 50:35]
      valid_7 <= 1'h0; // @[BPU.scala 52:16]
    end else if (io_wen) begin // @[BPU.scala 36:17]
      valid_7 <= _GEN_39;
    end
    if (reset) begin // @[BPU.scala 44:21]
      io_out_tag_REG <= 25'h0; // @[BPU.scala 44:21]
    end else if (3'h7 == io_index_r) begin // @[BPU.scala 44:21]
      io_out_tag_REG <= btb_entry_7_tag; // @[BPU.scala 44:21]
    end else if (3'h6 == io_index_r) begin // @[BPU.scala 44:21]
      io_out_tag_REG <= btb_entry_6_tag; // @[BPU.scala 44:21]
    end else if (3'h5 == io_index_r) begin // @[BPU.scala 44:21]
      io_out_tag_REG <= btb_entry_5_tag; // @[BPU.scala 44:21]
    end else begin
      io_out_tag_REG <= _GEN_84;
    end
    if (reset) begin // @[BPU.scala 45:24]
      io_out_offset_REG <= 2'h0; // @[BPU.scala 45:24]
    end else if (3'h7 == io_index_r) begin // @[BPU.scala 45:24]
      io_out_offset_REG <= btb_entry_7_offset; // @[BPU.scala 45:24]
    end else if (3'h6 == io_index_r) begin // @[BPU.scala 45:24]
      io_out_offset_REG <= btb_entry_6_offset; // @[BPU.scala 45:24]
    end else if (3'h5 == io_index_r) begin // @[BPU.scala 45:24]
      io_out_offset_REG <= btb_entry_5_offset; // @[BPU.scala 45:24]
    end else begin
      io_out_offset_REG <= _GEN_92;
    end
    if (reset) begin // @[BPU.scala 46:24]
      io_out_target_REG <= 32'h0; // @[BPU.scala 46:24]
    end else if (3'h7 == io_index_r) begin // @[BPU.scala 46:24]
      io_out_target_REG <= btb_entry_7_target; // @[BPU.scala 46:24]
    end else if (3'h6 == io_index_r) begin // @[BPU.scala 46:24]
      io_out_target_REG <= btb_entry_6_target; // @[BPU.scala 46:24]
    end else if (3'h5 == io_index_r) begin // @[BPU.scala 46:24]
      io_out_target_REG <= btb_entry_5_target; // @[BPU.scala 46:24]
    end else begin
      io_out_target_REG <= _GEN_100;
    end
    if (reset) begin // @[BPU.scala 47:26]
      io_out_btb_type_REG <= 2'h0; // @[BPU.scala 47:26]
    end else if (3'h7 == io_index_r) begin // @[BPU.scala 47:26]
      io_out_btb_type_REG <= btb_entry_7_btb_type; // @[BPU.scala 47:26]
    end else if (3'h6 == io_index_r) begin // @[BPU.scala 47:26]
      io_out_btb_type_REG <= btb_entry_6_btb_type; // @[BPU.scala 47:26]
    end else if (3'h5 == io_index_r) begin // @[BPU.scala 47:26]
      io_out_btb_type_REG <= btb_entry_5_btb_type; // @[BPU.scala 47:26]
    end else begin
      io_out_btb_type_REG <= _GEN_108;
    end
    if (reset) begin // @[BPU.scala 48:24]
      io_valid_r_REG <= 1'h0; // @[BPU.scala 48:24]
    end else if (3'h7 == io_index_r) begin // @[BPU.scala 48:24]
      io_valid_r_REG <= valid_7; // @[BPU.scala 48:24]
    end else if (3'h6 == io_index_r) begin // @[BPU.scala 48:24]
      io_valid_r_REG <= valid_6; // @[BPU.scala 48:24]
    end else if (3'h5 == io_index_r) begin // @[BPU.scala 48:24]
      io_valid_r_REG <= valid_5; // @[BPU.scala 48:24]
    end else begin
      io_valid_r_REG <= _GEN_116;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_entry_0_tag = _RAND_0[24:0];
  _RAND_1 = {1{`RANDOM}};
  btb_entry_0_offset = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  btb_entry_0_btb_type = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  btb_entry_0_target = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  btb_entry_1_tag = _RAND_4[24:0];
  _RAND_5 = {1{`RANDOM}};
  btb_entry_1_offset = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  btb_entry_1_btb_type = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  btb_entry_1_target = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  btb_entry_2_tag = _RAND_8[24:0];
  _RAND_9 = {1{`RANDOM}};
  btb_entry_2_offset = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  btb_entry_2_btb_type = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  btb_entry_2_target = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  btb_entry_3_tag = _RAND_12[24:0];
  _RAND_13 = {1{`RANDOM}};
  btb_entry_3_offset = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  btb_entry_3_btb_type = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  btb_entry_3_target = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  btb_entry_4_tag = _RAND_16[24:0];
  _RAND_17 = {1{`RANDOM}};
  btb_entry_4_offset = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  btb_entry_4_btb_type = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  btb_entry_4_target = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  btb_entry_5_tag = _RAND_20[24:0];
  _RAND_21 = {1{`RANDOM}};
  btb_entry_5_offset = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  btb_entry_5_btb_type = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  btb_entry_5_target = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  btb_entry_6_tag = _RAND_24[24:0];
  _RAND_25 = {1{`RANDOM}};
  btb_entry_6_offset = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  btb_entry_6_btb_type = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  btb_entry_6_target = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  btb_entry_7_tag = _RAND_28[24:0];
  _RAND_29 = {1{`RANDOM}};
  btb_entry_7_offset = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  btb_entry_7_btb_type = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  btb_entry_7_target = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  valid_0 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_1 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_3 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_4 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_5 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_6 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_7 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  io_out_tag_REG = _RAND_40[24:0];
  _RAND_41 = {1{`RANDOM}};
  io_out_offset_REG = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  io_out_target_REG = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  io_out_btb_type_REG = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  io_valid_r_REG = _RAND_44[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PHT(
  input        clock,
  input        reset,
  input        io_inc,
  input        io_dec,
  input  [3:0] io_index_w,
  input  [3:0] io_index_r,
  input        io_fence,
  output       io_br_taken
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pht_entry_0; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_1; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_2; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_3; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_4; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_5; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_6; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_7; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_8; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_9; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_10; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_11; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_12; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_13; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_14; // @[BPU.scala 69:26]
  reg [1:0] pht_entry_15; // @[BPU.scala 69:26]
  wire [1:0] _GEN_0 = reset | io_fence ? 2'h2 : pht_entry_0; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_1 = reset | io_fence ? 2'h2 : pht_entry_1; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_2 = reset | io_fence ? 2'h2 : pht_entry_2; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_3 = reset | io_fence ? 2'h2 : pht_entry_3; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_4 = reset | io_fence ? 2'h2 : pht_entry_4; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_5 = reset | io_fence ? 2'h2 : pht_entry_5; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_6 = reset | io_fence ? 2'h2 : pht_entry_6; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_7 = reset | io_fence ? 2'h2 : pht_entry_7; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_8 = reset | io_fence ? 2'h2 : pht_entry_8; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_9 = reset | io_fence ? 2'h2 : pht_entry_9; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_10 = reset | io_fence ? 2'h2 : pht_entry_10; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_11 = reset | io_fence ? 2'h2 : pht_entry_11; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_12 = reset | io_fence ? 2'h2 : pht_entry_12; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_13 = reset | io_fence ? 2'h2 : pht_entry_13; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_14 = reset | io_fence ? 2'h2 : pht_entry_14; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_15 = reset | io_fence ? 2'h2 : pht_entry_15; // @[BPU.scala 71:35 BPU.scala 73:20 BPU.scala 69:26]
  wire [1:0] _GEN_17 = 4'h1 == io_index_w ? pht_entry_1 : pht_entry_0; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_18 = 4'h2 == io_index_w ? pht_entry_2 : _GEN_17; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_19 = 4'h3 == io_index_w ? pht_entry_3 : _GEN_18; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_20 = 4'h4 == io_index_w ? pht_entry_4 : _GEN_19; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_21 = 4'h5 == io_index_w ? pht_entry_5 : _GEN_20; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_22 = 4'h6 == io_index_w ? pht_entry_6 : _GEN_21; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_23 = 4'h7 == io_index_w ? pht_entry_7 : _GEN_22; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_24 = 4'h8 == io_index_w ? pht_entry_8 : _GEN_23; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_25 = 4'h9 == io_index_w ? pht_entry_9 : _GEN_24; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_26 = 4'ha == io_index_w ? pht_entry_10 : _GEN_25; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_27 = 4'hb == io_index_w ? pht_entry_11 : _GEN_26; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_28 = 4'hc == io_index_w ? pht_entry_12 : _GEN_27; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_29 = 4'hd == io_index_w ? pht_entry_13 : _GEN_28; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_30 = 4'he == io_index_w ? pht_entry_14 : _GEN_29; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _GEN_31 = 4'hf == io_index_w ? pht_entry_15 : _GEN_30; // @[BPU.scala 78:50 BPU.scala 78:50]
  wire [1:0] _pht_entry_T_2 = _GEN_31 + 2'h1; // @[BPU.scala 78:91]
  wire [1:0] _pht_entry_T_6 = _GEN_31 - 2'h1; // @[BPU.scala 80:91]
  wire [1:0] _pht_entry_T_7 = _GEN_31 == 2'h0 ? 2'h0 : _pht_entry_T_6; // @[BPU.scala 80:30]
  wire [1:0] _GEN_97 = 4'h1 == io_index_r ? pht_entry_1 : pht_entry_0; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_98 = 4'h2 == io_index_r ? pht_entry_2 : _GEN_97; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_99 = 4'h3 == io_index_r ? pht_entry_3 : _GEN_98; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_100 = 4'h4 == io_index_r ? pht_entry_4 : _GEN_99; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_101 = 4'h5 == io_index_r ? pht_entry_5 : _GEN_100; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_102 = 4'h6 == io_index_r ? pht_entry_6 : _GEN_101; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_103 = 4'h7 == io_index_r ? pht_entry_7 : _GEN_102; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_104 = 4'h8 == io_index_r ? pht_entry_8 : _GEN_103; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_105 = 4'h9 == io_index_r ? pht_entry_9 : _GEN_104; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_106 = 4'ha == io_index_r ? pht_entry_10 : _GEN_105; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_107 = 4'hb == io_index_r ? pht_entry_11 : _GEN_106; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_108 = 4'hc == io_index_r ? pht_entry_12 : _GEN_107; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_109 = 4'hd == io_index_r ? pht_entry_13 : _GEN_108; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_110 = 4'he == io_index_r ? pht_entry_14 : _GEN_109; // @[BPU.scala 83:36 BPU.scala 83:36]
  wire [1:0] _GEN_111 = 4'hf == io_index_r ? pht_entry_15 : _GEN_110; // @[BPU.scala 83:36 BPU.scala 83:36]
  assign io_br_taken = _GEN_111[1]; // @[BPU.scala 83:36]
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_0 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h0 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_0 <= 2'h3;
        end else begin
          pht_entry_0 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_0 <= _GEN_0;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h0 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_0 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_0 <= _GEN_0;
      end
    end else begin
      pht_entry_0 <= _GEN_0;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_1 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h1 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_1 <= 2'h3;
        end else begin
          pht_entry_1 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_1 <= _GEN_1;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h1 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_1 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_1 <= _GEN_1;
      end
    end else begin
      pht_entry_1 <= _GEN_1;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_2 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h2 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_2 <= 2'h3;
        end else begin
          pht_entry_2 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_2 <= _GEN_2;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h2 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_2 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_2 <= _GEN_2;
      end
    end else begin
      pht_entry_2 <= _GEN_2;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_3 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h3 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_3 <= 2'h3;
        end else begin
          pht_entry_3 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_3 <= _GEN_3;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h3 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_3 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_3 <= _GEN_3;
      end
    end else begin
      pht_entry_3 <= _GEN_3;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_4 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h4 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_4 <= 2'h3;
        end else begin
          pht_entry_4 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_4 <= _GEN_4;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h4 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_4 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_4 <= _GEN_4;
      end
    end else begin
      pht_entry_4 <= _GEN_4;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_5 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h5 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_5 <= 2'h3;
        end else begin
          pht_entry_5 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_5 <= _GEN_5;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h5 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_5 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_5 <= _GEN_5;
      end
    end else begin
      pht_entry_5 <= _GEN_5;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_6 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h6 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_6 <= 2'h3;
        end else begin
          pht_entry_6 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_6 <= _GEN_6;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h6 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_6 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_6 <= _GEN_6;
      end
    end else begin
      pht_entry_6 <= _GEN_6;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_7 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h7 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_7 <= 2'h3;
        end else begin
          pht_entry_7 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_7 <= _GEN_7;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h7 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_7 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_7 <= _GEN_7;
      end
    end else begin
      pht_entry_7 <= _GEN_7;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_8 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h8 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_8 <= 2'h3;
        end else begin
          pht_entry_8 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_8 <= _GEN_8;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h8 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_8 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_8 <= _GEN_8;
      end
    end else begin
      pht_entry_8 <= _GEN_8;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_9 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'h9 == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_9 <= 2'h3;
        end else begin
          pht_entry_9 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_9 <= _GEN_9;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'h9 == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_9 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_9 <= _GEN_9;
      end
    end else begin
      pht_entry_9 <= _GEN_9;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_10 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'ha == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_10 <= 2'h3;
        end else begin
          pht_entry_10 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_10 <= _GEN_10;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'ha == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_10 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_10 <= _GEN_10;
      end
    end else begin
      pht_entry_10 <= _GEN_10;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_11 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'hb == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_11 <= 2'h3;
        end else begin
          pht_entry_11 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_11 <= _GEN_11;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'hb == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_11 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_11 <= _GEN_11;
      end
    end else begin
      pht_entry_11 <= _GEN_11;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_12 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'hc == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_12 <= 2'h3;
        end else begin
          pht_entry_12 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_12 <= _GEN_12;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'hc == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_12 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_12 <= _GEN_12;
      end
    end else begin
      pht_entry_12 <= _GEN_12;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_13 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'hd == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_13 <= 2'h3;
        end else begin
          pht_entry_13 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_13 <= _GEN_13;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'hd == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_13 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_13 <= _GEN_13;
      end
    end else begin
      pht_entry_13 <= _GEN_13;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_14 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'he == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_14 <= 2'h3;
        end else begin
          pht_entry_14 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_14 <= _GEN_14;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'he == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_14 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_14 <= _GEN_14;
      end
    end else begin
      pht_entry_14 <= _GEN_14;
    end
    if (reset) begin // @[BPU.scala 69:26]
      pht_entry_15 <= 2'h0; // @[BPU.scala 69:26]
    end else if (io_inc) begin // @[BPU.scala 77:17]
      if (4'hf == io_index_w) begin // @[BPU.scala 78:24]
        if (_GEN_31 == 2'h3) begin // @[BPU.scala 78:30]
          pht_entry_15 <= 2'h3;
        end else begin
          pht_entry_15 <= _pht_entry_T_2;
        end
      end else begin
        pht_entry_15 <= _GEN_15;
      end
    end else if (io_dec) begin // @[BPU.scala 79:24]
      if (4'hf == io_index_w) begin // @[BPU.scala 80:24]
        pht_entry_15 <= _pht_entry_T_7; // @[BPU.scala 80:24]
      end else begin
        pht_entry_15 <= _GEN_15;
      end
    end else begin
      pht_entry_15 <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pht_entry_0 = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  pht_entry_1 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  pht_entry_2 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  pht_entry_3 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  pht_entry_4 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  pht_entry_5 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  pht_entry_6 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  pht_entry_7 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  pht_entry_8 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  pht_entry_9 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  pht_entry_10 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  pht_entry_11 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  pht_entry_12 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  pht_entry_13 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  pht_entry_14 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  pht_entry_15 = _RAND_15[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RAS(
  input         clock,
  input         reset,
  input         io_call,
  input         io_ret,
  input  [2:0]  io_call_count,
  input  [2:0]  io_ret_count,
  input  [31:0] io_addr_w,
  output [31:0] io_addr_r,
  input         io_reflush,
  input         io_fence
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ras_entry_0; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_1; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_2; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_3; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_4; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_5; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_6; // @[BPU.scala 98:26]
  reg [31:0] ras_entry_7; // @[BPU.scala 98:26]
  wire  wrong_call = io_call_count > io_ret_count; // @[BPU.scala 103:31]
  wire [2:0] _wrong_count_T_1 = io_call_count - io_ret_count; // @[BPU.scala 106:48]
  wire [2:0] _wrong_count_T_3 = io_ret_count - io_call_count; // @[BPU.scala 106:77]
  wire [2:0] wrong_count = wrong_call ? _wrong_count_T_1 : _wrong_count_T_3; // @[BPU.scala 106:21]
  reg [2:0] ras_counter; // @[BPU.scala 108:28]
  wire [2:0] ras_counter_prev = ras_counter - 3'h1; // @[BPU.scala 115:35]
  wire [2:0] ras_counter_next = ras_counter + 3'h1; // @[BPU.scala 116:35]
  wire [31:0] _GEN_0 = reset | io_fence ? 32'h80000000 : ras_entry_0; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_1 = reset | io_fence ? 32'h80000000 : ras_entry_1; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_2 = reset | io_fence ? 32'h80000000 : ras_entry_2; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_3 = reset | io_fence ? 32'h80000000 : ras_entry_3; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_4 = reset | io_fence ? 32'h80000000 : ras_entry_4; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_5 = reset | io_fence ? 32'h80000000 : ras_entry_5; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_6 = reset | io_fence ? 32'h80000000 : ras_entry_6; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [31:0] _GEN_7 = reset | io_fence ? 32'h80000000 : ras_entry_7; // @[BPU.scala 120:35 BPU.scala 122:20 BPU.scala 98:26]
  wire [2:0] _GEN_8 = reset | io_fence ? 3'h0 : ras_counter; // @[BPU.scala 120:35 BPU.scala 124:17 BPU.scala 108:28]
  wire [2:0] _GEN_26 = io_ret ? ras_counter_prev : _GEN_8; // @[BPU.scala 132:24 BPU.scala 133:17]
  wire [2:0] _ras_counter_T_1 = ras_counter - wrong_count; // @[BPU.scala 137:32]
  wire [2:0] _ras_counter_T_3 = ras_counter + wrong_count; // @[BPU.scala 139:32]
  wire [31:0] _GEN_40 = 3'h1 == ras_counter_prev ? ras_entry_1 : ras_entry_0; // @[BPU.scala 142:13 BPU.scala 142:13]
  wire [31:0] _GEN_41 = 3'h2 == ras_counter_prev ? ras_entry_2 : _GEN_40; // @[BPU.scala 142:13 BPU.scala 142:13]
  wire [31:0] _GEN_42 = 3'h3 == ras_counter_prev ? ras_entry_3 : _GEN_41; // @[BPU.scala 142:13 BPU.scala 142:13]
  wire [31:0] _GEN_43 = 3'h4 == ras_counter_prev ? ras_entry_4 : _GEN_42; // @[BPU.scala 142:13 BPU.scala 142:13]
  wire [31:0] _GEN_44 = 3'h5 == ras_counter_prev ? ras_entry_5 : _GEN_43; // @[BPU.scala 142:13 BPU.scala 142:13]
  wire [31:0] _GEN_45 = 3'h6 == ras_counter_prev ? ras_entry_6 : _GEN_44; // @[BPU.scala 142:13 BPU.scala 142:13]
  assign io_addr_r = 3'h7 == ras_counter_prev ? ras_entry_7 : _GEN_45; // @[BPU.scala 142:13 BPU.scala 142:13]
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_0 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h0 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_0 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_0 <= _GEN_0;
      end
    end else begin
      ras_entry_0 <= _GEN_0;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_1 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h1 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_1 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_1 <= _GEN_1;
      end
    end else begin
      ras_entry_1 <= _GEN_1;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_2 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h2 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_2 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_2 <= _GEN_2;
      end
    end else begin
      ras_entry_2 <= _GEN_2;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_3 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h3 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_3 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_3 <= _GEN_3;
      end
    end else begin
      ras_entry_3 <= _GEN_3;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_4 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h4 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_4 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_4 <= _GEN_4;
      end
    end else begin
      ras_entry_4 <= _GEN_4;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_5 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h5 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_5 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_5 <= _GEN_5;
      end
    end else begin
      ras_entry_5 <= _GEN_5;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_6 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h6 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_6 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_6 <= _GEN_6;
      end
    end else begin
      ras_entry_6 <= _GEN_6;
    end
    if (reset) begin // @[BPU.scala 98:26]
      ras_entry_7 <= 32'h80000000; // @[BPU.scala 98:26]
    end else if (io_call) begin // @[BPU.scala 128:18]
      if (3'h7 == ras_counter) begin // @[BPU.scala 131:28]
        ras_entry_7 <= io_addr_w; // @[BPU.scala 131:28]
      end else begin
        ras_entry_7 <= _GEN_7;
      end
    end else begin
      ras_entry_7 <= _GEN_7;
    end
    if (reset) begin // @[BPU.scala 108:28]
      ras_counter <= 3'h0; // @[BPU.scala 108:28]
    end else if (io_reflush & wrong_call) begin // @[BPU.scala 136:35]
      ras_counter <= _ras_counter_T_1; // @[BPU.scala 137:17]
    end else if (io_reflush) begin // @[BPU.scala 138:28]
      ras_counter <= _ras_counter_T_3; // @[BPU.scala 139:17]
    end else if (io_call) begin // @[BPU.scala 128:18]
      ras_counter <= ras_counter_next; // @[BPU.scala 129:17]
    end else begin
      ras_counter <= _GEN_26;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ras_entry_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ras_entry_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ras_entry_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ras_entry_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  ras_entry_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  ras_entry_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  ras_entry_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ras_entry_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  ras_counter = _RAND_8[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BPU(
  input         clock,
  input         reset,
  input         io_ifu_valid,
  input  [31:0] io_ifu_pc,
  output        io_ifu_bp_ok,
  output        io_ifu_bp_taken,
  output [31:0] io_ifu_bp_target,
  output [1:0]  io_ifu_bp_offset,
  input         io_ifu_is_reflush,
  output [1:0]  io_ifu_bp_type,
  input  [2:0]  io_ifu_call_count,
  input  [2:0]  io_ifu_ret_count,
  input         io_exu_valid,
  input  [31:0] io_exu_pc,
  input         io_exu_bp_taken,
  input  [31:0] io_exu_bp_target,
  input  [1:0]  io_exu_bp_type,
  input         io_exu_bp_wrong,
  input         io_exu_fence,
  input  [2:0]  io_exu_call_count,
  input  [2:0]  io_exu_ret_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  wire  btb_0_clock; // @[BPU.scala 183:21]
  wire  btb_0_reset; // @[BPU.scala 183:21]
  wire  btb_0_io_wen; // @[BPU.scala 183:21]
  wire [2:0] btb_0_io_index_r; // @[BPU.scala 183:21]
  wire [2:0] btb_0_io_index_w; // @[BPU.scala 183:21]
  wire [24:0] btb_0_io_in_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_0_io_in_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_0_io_in_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_0_io_in_target; // @[BPU.scala 183:21]
  wire [24:0] btb_0_io_out_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_0_io_out_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_0_io_out_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_0_io_out_target; // @[BPU.scala 183:21]
  wire  btb_0_io_valid_r; // @[BPU.scala 183:21]
  wire  btb_0_io_fence; // @[BPU.scala 183:21]
  wire  btb_1_clock; // @[BPU.scala 183:21]
  wire  btb_1_reset; // @[BPU.scala 183:21]
  wire  btb_1_io_wen; // @[BPU.scala 183:21]
  wire [2:0] btb_1_io_index_r; // @[BPU.scala 183:21]
  wire [2:0] btb_1_io_index_w; // @[BPU.scala 183:21]
  wire [24:0] btb_1_io_in_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_1_io_in_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_1_io_in_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_1_io_in_target; // @[BPU.scala 183:21]
  wire [24:0] btb_1_io_out_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_1_io_out_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_1_io_out_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_1_io_out_target; // @[BPU.scala 183:21]
  wire  btb_1_io_valid_r; // @[BPU.scala 183:21]
  wire  btb_1_io_fence; // @[BPU.scala 183:21]
  wire  btb_2_clock; // @[BPU.scala 183:21]
  wire  btb_2_reset; // @[BPU.scala 183:21]
  wire  btb_2_io_wen; // @[BPU.scala 183:21]
  wire [2:0] btb_2_io_index_r; // @[BPU.scala 183:21]
  wire [2:0] btb_2_io_index_w; // @[BPU.scala 183:21]
  wire [24:0] btb_2_io_in_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_2_io_in_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_2_io_in_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_2_io_in_target; // @[BPU.scala 183:21]
  wire [24:0] btb_2_io_out_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_2_io_out_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_2_io_out_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_2_io_out_target; // @[BPU.scala 183:21]
  wire  btb_2_io_valid_r; // @[BPU.scala 183:21]
  wire  btb_2_io_fence; // @[BPU.scala 183:21]
  wire  btb_3_clock; // @[BPU.scala 183:21]
  wire  btb_3_reset; // @[BPU.scala 183:21]
  wire  btb_3_io_wen; // @[BPU.scala 183:21]
  wire [2:0] btb_3_io_index_r; // @[BPU.scala 183:21]
  wire [2:0] btb_3_io_index_w; // @[BPU.scala 183:21]
  wire [24:0] btb_3_io_in_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_3_io_in_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_3_io_in_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_3_io_in_target; // @[BPU.scala 183:21]
  wire [24:0] btb_3_io_out_tag; // @[BPU.scala 183:21]
  wire [1:0] btb_3_io_out_offset; // @[BPU.scala 183:21]
  wire [1:0] btb_3_io_out_btb_type; // @[BPU.scala 183:21]
  wire [31:0] btb_3_io_out_target; // @[BPU.scala 183:21]
  wire  btb_3_io_valid_r; // @[BPU.scala 183:21]
  wire  btb_3_io_fence; // @[BPU.scala 183:21]
  wire  pht_clock; // @[BPU.scala 195:19]
  wire  pht_reset; // @[BPU.scala 195:19]
  wire  pht_io_inc; // @[BPU.scala 195:19]
  wire  pht_io_dec; // @[BPU.scala 195:19]
  wire [3:0] pht_io_index_w; // @[BPU.scala 195:19]
  wire [3:0] pht_io_index_r; // @[BPU.scala 195:19]
  wire  pht_io_fence; // @[BPU.scala 195:19]
  wire  pht_io_br_taken; // @[BPU.scala 195:19]
  wire  ras_clock; // @[BPU.scala 202:19]
  wire  ras_reset; // @[BPU.scala 202:19]
  wire  ras_io_call; // @[BPU.scala 202:19]
  wire  ras_io_ret; // @[BPU.scala 202:19]
  wire [2:0] ras_io_call_count; // @[BPU.scala 202:19]
  wire [2:0] ras_io_ret_count; // @[BPU.scala 202:19]
  wire [31:0] ras_io_addr_w; // @[BPU.scala 202:19]
  wire [31:0] ras_io_addr_r; // @[BPU.scala 202:19]
  wire  ras_io_reflush; // @[BPU.scala 202:19]
  wire  ras_io_fence; // @[BPU.scala 202:19]
  reg [31:0] ifu_pc_reg; // @[BPU.scala 161:27]
  reg [31:0] exu_pc_reg; // @[BPU.scala 162:27]
  reg  exu_bp_taken_reg; // @[BPU.scala 163:33]
  reg [31:0] exu_bp_target_reg; // @[BPU.scala 164:34]
  reg [1:0] exu_bp_type_reg; // @[BPU.scala 165:32]
  reg  plru0_0; // @[BPU.scala 216:22]
  reg  plru0_1; // @[BPU.scala 216:22]
  reg  plru0_2; // @[BPU.scala 216:22]
  reg  plru0_3; // @[BPU.scala 216:22]
  reg  plru0_4; // @[BPU.scala 216:22]
  reg  plru0_5; // @[BPU.scala 216:22]
  reg  plru0_6; // @[BPU.scala 216:22]
  reg  plru0_7; // @[BPU.scala 216:22]
  reg  plru1_0; // @[BPU.scala 217:22]
  reg  plru1_1; // @[BPU.scala 217:22]
  reg  plru1_2; // @[BPU.scala 217:22]
  reg  plru1_3; // @[BPU.scala 217:22]
  reg  plru1_4; // @[BPU.scala 217:22]
  reg  plru1_5; // @[BPU.scala 217:22]
  reg  plru1_6; // @[BPU.scala 217:22]
  reg  plru1_7; // @[BPU.scala 217:22]
  reg  plru2_0; // @[BPU.scala 218:22]
  reg  plru2_1; // @[BPU.scala 218:22]
  reg  plru2_2; // @[BPU.scala 218:22]
  reg  plru2_3; // @[BPU.scala 218:22]
  reg  plru2_4; // @[BPU.scala 218:22]
  reg  plru2_5; // @[BPU.scala 218:22]
  reg  plru2_6; // @[BPU.scala 218:22]
  reg  plru2_7; // @[BPU.scala 218:22]
  reg [1:0] ifu_state; // @[BPU.scala 234:26]
  reg [1:0] exu_state; // @[BPU.scala 235:26]
  wire [24:0] tag_0 = btb_0_io_out_tag;
  wire  valid_0 = btb_0_io_valid_r;
  wire  ifu_hit_0 = tag_0 == ifu_pc_reg[31:7] & valid_0; // @[BPU.scala 238:42]
  wire [24:0] tag_1 = btb_1_io_out_tag;
  wire  valid_1 = btb_1_io_valid_r;
  wire  ifu_hit_1 = tag_1 == ifu_pc_reg[31:7] & valid_1; // @[BPU.scala 238:42]
  wire [24:0] tag_2 = btb_2_io_out_tag;
  wire  valid_2 = btb_2_io_valid_r;
  wire  ifu_hit_2 = tag_2 == ifu_pc_reg[31:7] & valid_2; // @[BPU.scala 238:42]
  wire [24:0] tag_3 = btb_3_io_out_tag;
  wire  valid_3 = btb_3_io_valid_r;
  wire  ifu_hit_3 = tag_3 == ifu_pc_reg[31:7] & valid_3; // @[BPU.scala 238:42]
  wire [3:0] _ifu_btb_hit_T = {ifu_hit_0,ifu_hit_1,ifu_hit_2,ifu_hit_3}; // @[Cat.scala 30:58]
  wire  ifu_btb_hit = |_ifu_btb_hit_T; // @[BPU.scala 240:31]
  wire  exu_hit_0 = tag_0 == exu_pc_reg[31:7] & valid_0; // @[BPU.scala 243:42]
  wire  exu_hit_1 = tag_1 == exu_pc_reg[31:7] & valid_1; // @[BPU.scala 243:42]
  wire  exu_hit_2 = tag_2 == exu_pc_reg[31:7] & valid_2; // @[BPU.scala 243:42]
  wire  exu_hit_3 = tag_3 == exu_pc_reg[31:7] & valid_3; // @[BPU.scala 243:42]
  wire [3:0] _exu_btb_hit_T = {exu_hit_0,exu_hit_1,exu_hit_2,exu_hit_3}; // @[Cat.scala 30:58]
  wire  exu_btb_hit = |_exu_btb_hit_T; // @[BPU.scala 245:31]
  wire  _GEN_7 = 3'h0 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_0; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_8 = 3'h1 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_1; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_9 = 3'h2 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_2; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_10 = 3'h3 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_3; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_11 = 3'h4 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_4; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_12 = 3'h5 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_5; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_13 = 3'h6 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_6; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_14 = 3'h7 == exu_pc_reg[6:4] ? exu_hit_0 | exu_hit_1 : plru0_7; // @[BPU.scala 248:38 BPU.scala 248:38 BPU.scala 216:22]
  wire  _GEN_583 = 3'h0 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_15 = 3'h0 == exu_pc_reg[6:4] | plru1_0; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_584 = 3'h1 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_16 = 3'h1 == exu_pc_reg[6:4] | plru1_1; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_585 = 3'h2 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_17 = 3'h2 == exu_pc_reg[6:4] | plru1_2; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_586 = 3'h3 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_18 = 3'h3 == exu_pc_reg[6:4] | plru1_3; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_587 = 3'h4 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_19 = 3'h4 == exu_pc_reg[6:4] | plru1_4; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_588 = 3'h5 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_20 = 3'h5 == exu_pc_reg[6:4] | plru1_5; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_589 = 3'h6 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_21 = 3'h6 == exu_pc_reg[6:4] | plru1_6; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_590 = 3'h7 == exu_pc_reg[6:4]; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_22 = 3'h7 == exu_pc_reg[6:4] | plru1_7; // @[BPU.scala 250:40 BPU.scala 250:40 BPU.scala 217:22]
  wire  _GEN_23 = 3'h0 == exu_pc_reg[6:4] ? 1'h0 : plru1_0; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_24 = 3'h1 == exu_pc_reg[6:4] ? 1'h0 : plru1_1; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_25 = 3'h2 == exu_pc_reg[6:4] ? 1'h0 : plru1_2; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_26 = 3'h3 == exu_pc_reg[6:4] ? 1'h0 : plru1_3; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_27 = 3'h4 == exu_pc_reg[6:4] ? 1'h0 : plru1_4; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_28 = 3'h5 == exu_pc_reg[6:4] ? 1'h0 : plru1_5; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_29 = 3'h6 == exu_pc_reg[6:4] ? 1'h0 : plru1_6; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_30 = 3'h7 == exu_pc_reg[6:4] ? 1'h0 : plru1_7; // @[BPU.scala 252:40 BPU.scala 252:40 BPU.scala 217:22]
  wire  _GEN_31 = _GEN_583 | plru2_0; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_32 = _GEN_584 | plru2_1; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_33 = _GEN_585 | plru2_2; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_34 = _GEN_586 | plru2_3; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_35 = _GEN_587 | plru2_4; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_36 = _GEN_588 | plru2_5; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_37 = _GEN_589 | plru2_6; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_38 = _GEN_590 | plru2_7; // @[BPU.scala 254:40 BPU.scala 254:40 BPU.scala 218:22]
  wire  _GEN_39 = 3'h0 == exu_pc_reg[6:4] ? 1'h0 : plru2_0; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_40 = 3'h1 == exu_pc_reg[6:4] ? 1'h0 : plru2_1; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_41 = 3'h2 == exu_pc_reg[6:4] ? 1'h0 : plru2_2; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_42 = 3'h3 == exu_pc_reg[6:4] ? 1'h0 : plru2_3; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_43 = 3'h4 == exu_pc_reg[6:4] ? 1'h0 : plru2_4; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_44 = 3'h5 == exu_pc_reg[6:4] ? 1'h0 : plru2_5; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_45 = 3'h6 == exu_pc_reg[6:4] ? 1'h0 : plru2_6; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_46 = 3'h7 == exu_pc_reg[6:4] ? 1'h0 : plru2_7; // @[BPU.scala 256:40 BPU.scala 256:40 BPU.scala 218:22]
  wire  _GEN_47 = exu_hit_3 ? _GEN_39 : plru2_0; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_48 = exu_hit_3 ? _GEN_40 : plru2_1; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_49 = exu_hit_3 ? _GEN_41 : plru2_2; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_50 = exu_hit_3 ? _GEN_42 : plru2_3; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_51 = exu_hit_3 ? _GEN_43 : plru2_4; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_52 = exu_hit_3 ? _GEN_44 : plru2_5; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_53 = exu_hit_3 ? _GEN_45 : plru2_6; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_54 = exu_hit_3 ? _GEN_46 : plru2_7; // @[BPU.scala 255:30 BPU.scala 218:22]
  wire  _GEN_55 = exu_hit_2 ? _GEN_31 : _GEN_47; // @[BPU.scala 253:30]
  wire  _GEN_56 = exu_hit_2 ? _GEN_32 : _GEN_48; // @[BPU.scala 253:30]
  wire  _GEN_57 = exu_hit_2 ? _GEN_33 : _GEN_49; // @[BPU.scala 253:30]
  wire  _GEN_58 = exu_hit_2 ? _GEN_34 : _GEN_50; // @[BPU.scala 253:30]
  wire  _GEN_59 = exu_hit_2 ? _GEN_35 : _GEN_51; // @[BPU.scala 253:30]
  wire  _GEN_60 = exu_hit_2 ? _GEN_36 : _GEN_52; // @[BPU.scala 253:30]
  wire  _GEN_61 = exu_hit_2 ? _GEN_37 : _GEN_53; // @[BPU.scala 253:30]
  wire  _GEN_62 = exu_hit_2 ? _GEN_38 : _GEN_54; // @[BPU.scala 253:30]
  wire  _GEN_63 = exu_hit_1 ? _GEN_23 : plru1_0; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_64 = exu_hit_1 ? _GEN_24 : plru1_1; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_65 = exu_hit_1 ? _GEN_25 : plru1_2; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_66 = exu_hit_1 ? _GEN_26 : plru1_3; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_67 = exu_hit_1 ? _GEN_27 : plru1_4; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_68 = exu_hit_1 ? _GEN_28 : plru1_5; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_69 = exu_hit_1 ? _GEN_29 : plru1_6; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_70 = exu_hit_1 ? _GEN_30 : plru1_7; // @[BPU.scala 251:30 BPU.scala 217:22]
  wire  _GEN_71 = exu_hit_1 ? plru2_0 : _GEN_55; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_72 = exu_hit_1 ? plru2_1 : _GEN_56; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_73 = exu_hit_1 ? plru2_2 : _GEN_57; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_74 = exu_hit_1 ? plru2_3 : _GEN_58; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_75 = exu_hit_1 ? plru2_4 : _GEN_59; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_76 = exu_hit_1 ? plru2_5 : _GEN_60; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_77 = exu_hit_1 ? plru2_6 : _GEN_61; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_78 = exu_hit_1 ? plru2_7 : _GEN_62; // @[BPU.scala 251:30 BPU.scala 218:22]
  wire  _GEN_79 = exu_hit_0 ? _GEN_15 : _GEN_63; // @[BPU.scala 249:23]
  wire  _GEN_80 = exu_hit_0 ? _GEN_16 : _GEN_64; // @[BPU.scala 249:23]
  wire  _GEN_81 = exu_hit_0 ? _GEN_17 : _GEN_65; // @[BPU.scala 249:23]
  wire  _GEN_82 = exu_hit_0 ? _GEN_18 : _GEN_66; // @[BPU.scala 249:23]
  wire  _GEN_83 = exu_hit_0 ? _GEN_19 : _GEN_67; // @[BPU.scala 249:23]
  wire  _GEN_84 = exu_hit_0 ? _GEN_20 : _GEN_68; // @[BPU.scala 249:23]
  wire  _GEN_85 = exu_hit_0 ? _GEN_21 : _GEN_69; // @[BPU.scala 249:23]
  wire  _GEN_86 = exu_hit_0 ? _GEN_22 : _GEN_70; // @[BPU.scala 249:23]
  wire  _GEN_87 = exu_hit_0 ? plru2_0 : _GEN_71; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_88 = exu_hit_0 ? plru2_1 : _GEN_72; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_89 = exu_hit_0 ? plru2_2 : _GEN_73; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_90 = exu_hit_0 ? plru2_3 : _GEN_74; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_91 = exu_hit_0 ? plru2_4 : _GEN_75; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_92 = exu_hit_0 ? plru2_5 : _GEN_76; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_93 = exu_hit_0 ? plru2_6 : _GEN_77; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_94 = exu_hit_0 ? plru2_7 : _GEN_78; // @[BPU.scala 249:23 BPU.scala 218:22]
  wire  _GEN_95 = exu_state == 2'h1 & exu_btb_hit ? _GEN_7 : plru0_0; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_96 = exu_state == 2'h1 & exu_btb_hit ? _GEN_8 : plru0_1; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_97 = exu_state == 2'h1 & exu_btb_hit ? _GEN_9 : plru0_2; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_98 = exu_state == 2'h1 & exu_btb_hit ? _GEN_10 : plru0_3; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_99 = exu_state == 2'h1 & exu_btb_hit ? _GEN_11 : plru0_4; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_100 = exu_state == 2'h1 & exu_btb_hit ? _GEN_12 : plru0_5; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_101 = exu_state == 2'h1 & exu_btb_hit ? _GEN_13 : plru0_6; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_102 = exu_state == 2'h1 & exu_btb_hit ? _GEN_14 : plru0_7; // @[BPU.scala 247:55 BPU.scala 216:22]
  wire  _GEN_103 = exu_state == 2'h1 & exu_btb_hit ? _GEN_79 : plru1_0; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_104 = exu_state == 2'h1 & exu_btb_hit ? _GEN_80 : plru1_1; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_105 = exu_state == 2'h1 & exu_btb_hit ? _GEN_81 : plru1_2; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_106 = exu_state == 2'h1 & exu_btb_hit ? _GEN_82 : plru1_3; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_107 = exu_state == 2'h1 & exu_btb_hit ? _GEN_83 : plru1_4; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_108 = exu_state == 2'h1 & exu_btb_hit ? _GEN_84 : plru1_5; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_109 = exu_state == 2'h1 & exu_btb_hit ? _GEN_85 : plru1_6; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_110 = exu_state == 2'h1 & exu_btb_hit ? _GEN_86 : plru1_7; // @[BPU.scala 247:55 BPU.scala 217:22]
  wire  _GEN_111 = exu_state == 2'h1 & exu_btb_hit ? _GEN_87 : plru2_0; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_112 = exu_state == 2'h1 & exu_btb_hit ? _GEN_88 : plru2_1; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_113 = exu_state == 2'h1 & exu_btb_hit ? _GEN_89 : plru2_2; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_114 = exu_state == 2'h1 & exu_btb_hit ? _GEN_90 : plru2_3; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_115 = exu_state == 2'h1 & exu_btb_hit ? _GEN_91 : plru2_4; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_116 = exu_state == 2'h1 & exu_btb_hit ? _GEN_92 : plru2_5; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_117 = exu_state == 2'h1 & exu_btb_hit ? _GEN_93 : plru2_6; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_118 = exu_state == 2'h1 & exu_btb_hit ? _GEN_94 : plru2_7; // @[BPU.scala 247:55 BPU.scala 218:22]
  wire  _GEN_599 = 3'h0 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_127 = 3'h0 == ifu_pc_reg[6:4] | _GEN_103; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_600 = 3'h1 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_128 = 3'h1 == ifu_pc_reg[6:4] | _GEN_104; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_601 = 3'h2 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_129 = 3'h2 == ifu_pc_reg[6:4] | _GEN_105; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_602 = 3'h3 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_130 = 3'h3 == ifu_pc_reg[6:4] | _GEN_106; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_603 = 3'h4 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_131 = 3'h4 == ifu_pc_reg[6:4] | _GEN_107; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_604 = 3'h5 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_132 = 3'h5 == ifu_pc_reg[6:4] | _GEN_108; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_605 = 3'h6 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_133 = 3'h6 == ifu_pc_reg[6:4] | _GEN_109; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_606 = 3'h7 == ifu_pc_reg[6:4]; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_134 = 3'h7 == ifu_pc_reg[6:4] | _GEN_110; // @[BPU.scala 263:40 BPU.scala 263:40]
  wire  _GEN_135 = 3'h0 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_103; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_136 = 3'h1 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_104; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_137 = 3'h2 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_105; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_138 = 3'h3 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_106; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_139 = 3'h4 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_107; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_140 = 3'h5 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_108; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_141 = 3'h6 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_109; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_142 = 3'h7 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_110; // @[BPU.scala 265:40 BPU.scala 265:40]
  wire  _GEN_143 = _GEN_599 | _GEN_111; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_144 = _GEN_600 | _GEN_112; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_145 = _GEN_601 | _GEN_113; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_146 = _GEN_602 | _GEN_114; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_147 = _GEN_603 | _GEN_115; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_148 = _GEN_604 | _GEN_116; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_149 = _GEN_605 | _GEN_117; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_150 = _GEN_606 | _GEN_118; // @[BPU.scala 267:40 BPU.scala 267:40]
  wire  _GEN_151 = 3'h0 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_111; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_152 = 3'h1 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_112; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_153 = 3'h2 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_113; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_154 = 3'h3 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_114; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_155 = 3'h4 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_115; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_156 = 3'h5 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_116; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_157 = 3'h6 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_117; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_158 = 3'h7 == ifu_pc_reg[6:4] ? 1'h0 : _GEN_118; // @[BPU.scala 269:40 BPU.scala 269:40]
  wire  _GEN_159 = ifu_hit_3 ? _GEN_151 : _GEN_111; // @[BPU.scala 268:30]
  wire  _GEN_160 = ifu_hit_3 ? _GEN_152 : _GEN_112; // @[BPU.scala 268:30]
  wire  _GEN_161 = ifu_hit_3 ? _GEN_153 : _GEN_113; // @[BPU.scala 268:30]
  wire  _GEN_162 = ifu_hit_3 ? _GEN_154 : _GEN_114; // @[BPU.scala 268:30]
  wire  _GEN_163 = ifu_hit_3 ? _GEN_155 : _GEN_115; // @[BPU.scala 268:30]
  wire  _GEN_164 = ifu_hit_3 ? _GEN_156 : _GEN_116; // @[BPU.scala 268:30]
  wire  _GEN_165 = ifu_hit_3 ? _GEN_157 : _GEN_117; // @[BPU.scala 268:30]
  wire  _GEN_166 = ifu_hit_3 ? _GEN_158 : _GEN_118; // @[BPU.scala 268:30]
  wire  _GEN_167 = ifu_hit_2 ? _GEN_143 : _GEN_159; // @[BPU.scala 266:30]
  wire  _GEN_168 = ifu_hit_2 ? _GEN_144 : _GEN_160; // @[BPU.scala 266:30]
  wire  _GEN_169 = ifu_hit_2 ? _GEN_145 : _GEN_161; // @[BPU.scala 266:30]
  wire  _GEN_170 = ifu_hit_2 ? _GEN_146 : _GEN_162; // @[BPU.scala 266:30]
  wire  _GEN_171 = ifu_hit_2 ? _GEN_147 : _GEN_163; // @[BPU.scala 266:30]
  wire  _GEN_172 = ifu_hit_2 ? _GEN_148 : _GEN_164; // @[BPU.scala 266:30]
  wire  _GEN_173 = ifu_hit_2 ? _GEN_149 : _GEN_165; // @[BPU.scala 266:30]
  wire  _GEN_174 = ifu_hit_2 ? _GEN_150 : _GEN_166; // @[BPU.scala 266:30]
  wire  _GEN_232 = 3'h1 == exu_pc_reg[6:4] ? plru0_1 : plru0_0; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_233 = 3'h2 == exu_pc_reg[6:4] ? plru0_2 : _GEN_232; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_234 = 3'h3 == exu_pc_reg[6:4] ? plru0_3 : _GEN_233; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_235 = 3'h4 == exu_pc_reg[6:4] ? plru0_4 : _GEN_234; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_236 = 3'h5 == exu_pc_reg[6:4] ? plru0_5 : _GEN_235; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_237 = 3'h6 == exu_pc_reg[6:4] ? plru0_6 : _GEN_236; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_238 = 3'h7 == exu_pc_reg[6:4] ? plru0_7 : _GEN_237; // @[BPU.scala 274:42 BPU.scala 274:42]
  wire  _GEN_240 = 3'h1 == exu_pc_reg[6:4] ? plru1_1 : plru1_0; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_241 = 3'h2 == exu_pc_reg[6:4] ? plru1_2 : _GEN_240; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_242 = 3'h3 == exu_pc_reg[6:4] ? plru1_3 : _GEN_241; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_243 = 3'h4 == exu_pc_reg[6:4] ? plru1_4 : _GEN_242; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_244 = 3'h5 == exu_pc_reg[6:4] ? plru1_5 : _GEN_243; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_245 = 3'h6 == exu_pc_reg[6:4] ? plru1_6 : _GEN_244; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_246 = 3'h7 == exu_pc_reg[6:4] ? plru1_7 : _GEN_245; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_248 = 3'h1 == exu_pc_reg[6:4] ? plru2_1 : plru2_0; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_249 = 3'h2 == exu_pc_reg[6:4] ? plru2_2 : _GEN_248; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_250 = 3'h3 == exu_pc_reg[6:4] ? plru2_3 : _GEN_249; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_251 = 3'h4 == exu_pc_reg[6:4] ? plru2_4 : _GEN_250; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_252 = 3'h5 == exu_pc_reg[6:4] ? plru2_5 : _GEN_251; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_253 = 3'h6 == exu_pc_reg[6:4] ? plru2_6 : _GEN_252; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  _GEN_254 = 3'h7 == exu_pc_reg[6:4] ? plru2_7 : _GEN_253; // @[BPU.scala 274:8 BPU.scala 274:8]
  wire  replace_way_lo = ~_GEN_238 ? _GEN_246 : _GEN_254; // @[BPU.scala 274:8]
  wire [1:0] replace_way = {_GEN_238,replace_way_lo}; // @[Cat.scala 30:58]
  wire  _T_14 = 2'h0 == exu_state; // @[Conditional.scala 37:30]
  wire  _T_15 = io_exu_valid & io_exu_bp_wrong; // @[BPU.scala 284:23]
  wire [2:0] _GEN_265 = io_exu_valid & io_exu_bp_wrong ? io_exu_pc[6:4] : 3'h0; // @[BPU.scala 284:40 BPU.scala 287:29 BPU.scala 189:18]
  wire  _T_16 = 2'h1 == exu_state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_269 = exu_bp_type_reg == 2'h2 ? exu_pc_reg[7:4] : 4'h0; // @[BPU.scala 295:47 BPU.scala 296:26 BPU.scala 198:18]
  wire  _GEN_270 = exu_bp_type_reg == 2'h2 & exu_bp_taken_reg; // @[BPU.scala 295:47 BPU.scala 297:22 BPU.scala 196:14]
  wire  _GEN_271 = exu_bp_type_reg == 2'h2 & ~exu_bp_taken_reg; // @[BPU.scala 295:47 BPU.scala 298:22 BPU.scala 197:14]
  wire  _T_18 = replace_way == 2'h0; // @[BPU.scala 305:29]
  wire [2:0] _GEN_273 = replace_way == 2'h0 ? exu_pc_reg[6:4] : 3'h0; // @[BPU.scala 305:38 BPU.scala 307:31 BPU.scala 190:18]
  wire [24:0] _GEN_274 = replace_way == 2'h0 ? exu_pc_reg[31:7] : 25'h0; // @[BPU.scala 305:38 BPU.scala 308:30 BPU.scala 191:13]
  wire [1:0] _GEN_275 = replace_way == 2'h0 ? exu_pc_reg[3:2] : 2'h0; // @[BPU.scala 305:38 BPU.scala 309:33 BPU.scala 191:13]
  wire [1:0] _GEN_276 = replace_way == 2'h0 ? exu_bp_type_reg : 2'h0; // @[BPU.scala 305:38 BPU.scala 310:35 BPU.scala 191:13]
  wire [31:0] _GEN_277 = replace_way == 2'h0 ? exu_bp_target_reg : 32'h0; // @[BPU.scala 305:38 BPU.scala 311:33 BPU.scala 191:13]
  wire  _T_19 = replace_way == 2'h1; // @[BPU.scala 305:29]
  wire [2:0] _GEN_279 = replace_way == 2'h1 ? exu_pc_reg[6:4] : 3'h0; // @[BPU.scala 305:38 BPU.scala 307:31 BPU.scala 190:18]
  wire [24:0] _GEN_280 = replace_way == 2'h1 ? exu_pc_reg[31:7] : 25'h0; // @[BPU.scala 305:38 BPU.scala 308:30 BPU.scala 191:13]
  wire [1:0] _GEN_281 = replace_way == 2'h1 ? exu_pc_reg[3:2] : 2'h0; // @[BPU.scala 305:38 BPU.scala 309:33 BPU.scala 191:13]
  wire [1:0] _GEN_282 = replace_way == 2'h1 ? exu_bp_type_reg : 2'h0; // @[BPU.scala 305:38 BPU.scala 310:35 BPU.scala 191:13]
  wire [31:0] _GEN_283 = replace_way == 2'h1 ? exu_bp_target_reg : 32'h0; // @[BPU.scala 305:38 BPU.scala 311:33 BPU.scala 191:13]
  wire  _T_20 = replace_way == 2'h2; // @[BPU.scala 305:29]
  wire [2:0] _GEN_285 = replace_way == 2'h2 ? exu_pc_reg[6:4] : 3'h0; // @[BPU.scala 305:38 BPU.scala 307:31 BPU.scala 190:18]
  wire [24:0] _GEN_286 = replace_way == 2'h2 ? exu_pc_reg[31:7] : 25'h0; // @[BPU.scala 305:38 BPU.scala 308:30 BPU.scala 191:13]
  wire [1:0] _GEN_287 = replace_way == 2'h2 ? exu_pc_reg[3:2] : 2'h0; // @[BPU.scala 305:38 BPU.scala 309:33 BPU.scala 191:13]
  wire [1:0] _GEN_288 = replace_way == 2'h2 ? exu_bp_type_reg : 2'h0; // @[BPU.scala 305:38 BPU.scala 310:35 BPU.scala 191:13]
  wire [31:0] _GEN_289 = replace_way == 2'h2 ? exu_bp_target_reg : 32'h0; // @[BPU.scala 305:38 BPU.scala 311:33 BPU.scala 191:13]
  wire  _T_21 = replace_way == 2'h3; // @[BPU.scala 305:29]
  wire [2:0] _GEN_291 = replace_way == 2'h3 ? exu_pc_reg[6:4] : 3'h0; // @[BPU.scala 305:38 BPU.scala 307:31 BPU.scala 190:18]
  wire [24:0] _GEN_292 = replace_way == 2'h3 ? exu_pc_reg[31:7] : 25'h0; // @[BPU.scala 305:38 BPU.scala 308:30 BPU.scala 191:13]
  wire [1:0] _GEN_293 = replace_way == 2'h3 ? exu_pc_reg[3:2] : 2'h0; // @[BPU.scala 305:38 BPU.scala 309:33 BPU.scala 191:13]
  wire [1:0] _GEN_294 = replace_way == 2'h3 ? exu_bp_type_reg : 2'h0; // @[BPU.scala 305:38 BPU.scala 310:35 BPU.scala 191:13]
  wire [31:0] _GEN_295 = replace_way == 2'h3 ? exu_bp_target_reg : 32'h0; // @[BPU.scala 305:38 BPU.scala 311:33 BPU.scala 191:13]
  wire [3:0] _GEN_299 = exu_btb_hit ? _GEN_269 : _GEN_269; // @[BPU.scala 294:26]
  wire  _GEN_300 = exu_btb_hit ? _GEN_270 : _GEN_270; // @[BPU.scala 294:26]
  wire  _GEN_301 = exu_btb_hit ? _GEN_271 : _GEN_271; // @[BPU.scala 294:26]
  wire  _GEN_303 = exu_btb_hit ? 1'h0 : _T_18; // @[BPU.scala 294:26 BPU.scala 188:14]
  wire [2:0] _GEN_304 = exu_btb_hit ? 3'h0 : _GEN_273; // @[BPU.scala 294:26 BPU.scala 190:18]
  wire [24:0] _GEN_305 = exu_btb_hit ? 25'h0 : _GEN_274; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_306 = exu_btb_hit ? 2'h0 : _GEN_275; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_307 = exu_btb_hit ? 2'h0 : _GEN_276; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [31:0] _GEN_308 = exu_btb_hit ? 32'h0 : _GEN_277; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire  _GEN_309 = exu_btb_hit ? 1'h0 : _T_19; // @[BPU.scala 294:26 BPU.scala 188:14]
  wire [2:0] _GEN_310 = exu_btb_hit ? 3'h0 : _GEN_279; // @[BPU.scala 294:26 BPU.scala 190:18]
  wire [24:0] _GEN_311 = exu_btb_hit ? 25'h0 : _GEN_280; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_312 = exu_btb_hit ? 2'h0 : _GEN_281; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_313 = exu_btb_hit ? 2'h0 : _GEN_282; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [31:0] _GEN_314 = exu_btb_hit ? 32'h0 : _GEN_283; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire  _GEN_315 = exu_btb_hit ? 1'h0 : _T_20; // @[BPU.scala 294:26 BPU.scala 188:14]
  wire [2:0] _GEN_316 = exu_btb_hit ? 3'h0 : _GEN_285; // @[BPU.scala 294:26 BPU.scala 190:18]
  wire [24:0] _GEN_317 = exu_btb_hit ? 25'h0 : _GEN_286; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_318 = exu_btb_hit ? 2'h0 : _GEN_287; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_319 = exu_btb_hit ? 2'h0 : _GEN_288; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [31:0] _GEN_320 = exu_btb_hit ? 32'h0 : _GEN_289; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire  _GEN_321 = exu_btb_hit ? 1'h0 : _T_21; // @[BPU.scala 294:26 BPU.scala 188:14]
  wire [2:0] _GEN_322 = exu_btb_hit ? 3'h0 : _GEN_291; // @[BPU.scala 294:26 BPU.scala 190:18]
  wire [24:0] _GEN_323 = exu_btb_hit ? 25'h0 : _GEN_292; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_324 = exu_btb_hit ? 2'h0 : _GEN_293; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [1:0] _GEN_325 = exu_btb_hit ? 2'h0 : _GEN_294; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire [31:0] _GEN_326 = exu_btb_hit ? 32'h0 : _GEN_295; // @[BPU.scala 294:26 BPU.scala 191:13]
  wire  _T_23 = exu_bp_type_reg == 2'h0; // @[BPU.scala 324:29]
  wire [31:0] _ras_io_addr_w_T_1 = exu_pc_reg + 32'h4; // @[BPU.scala 326:37]
  wire  _T_24 = exu_bp_type_reg == 2'h1; // @[BPU.scala 327:36]
  wire [31:0] _GEN_329 = exu_bp_type_reg == 2'h0 ? _ras_io_addr_w_T_1 : 32'h0; // @[BPU.scala 324:43 BPU.scala 326:23 BPU.scala 205:17]
  wire  _GEN_330 = exu_bp_type_reg == 2'h0 ? 1'h0 : _T_24; // @[BPU.scala 324:43 BPU.scala 204:14]
  wire  _T_25 = 2'h2 == exu_state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_334 = io_exu_valid ? 2'h2 : 2'h0; // @[BPU.scala 344:31 BPU.scala 345:19 BPU.scala 347:19]
  wire [1:0] _GEN_335 = _T_15 ? 2'h1 : _GEN_334; // @[BPU.scala 339:40 BPU.scala 340:19]
  wire [3:0] _GEN_340 = _T_25 ? _GEN_269 : 4'h0; // @[Conditional.scala 39:67 BPU.scala 198:18]
  wire  _GEN_341 = _T_25 & _GEN_270; // @[Conditional.scala 39:67 BPU.scala 196:14]
  wire  _GEN_342 = _T_25 & _GEN_271; // @[Conditional.scala 39:67 BPU.scala 197:14]
  wire [2:0] _GEN_344 = _T_25 ? _GEN_265 : 3'h0; // @[Conditional.scala 39:67 BPU.scala 189:18]
  wire [3:0] _GEN_348 = _T_16 ? _GEN_299 : _GEN_340; // @[Conditional.scala 39:67]
  wire  _GEN_349 = _T_16 ? _GEN_300 : _GEN_341; // @[Conditional.scala 39:67]
  wire  _GEN_350 = _T_16 ? _GEN_301 : _GEN_342; // @[Conditional.scala 39:67]
  wire  _GEN_352 = _T_16 & _GEN_303; // @[Conditional.scala 39:67 BPU.scala 188:14]
  wire [2:0] _GEN_353 = _T_16 ? _GEN_304 : 3'h0; // @[Conditional.scala 39:67 BPU.scala 190:18]
  wire [24:0] _GEN_354 = _T_16 ? _GEN_305 : 25'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_355 = _T_16 ? _GEN_306 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_356 = _T_16 ? _GEN_307 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [31:0] _GEN_357 = _T_16 ? _GEN_308 : 32'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire  _GEN_358 = _T_16 & _GEN_309; // @[Conditional.scala 39:67 BPU.scala 188:14]
  wire [2:0] _GEN_359 = _T_16 ? _GEN_310 : 3'h0; // @[Conditional.scala 39:67 BPU.scala 190:18]
  wire [24:0] _GEN_360 = _T_16 ? _GEN_311 : 25'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_361 = _T_16 ? _GEN_312 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_362 = _T_16 ? _GEN_313 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [31:0] _GEN_363 = _T_16 ? _GEN_314 : 32'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire  _GEN_364 = _T_16 & _GEN_315; // @[Conditional.scala 39:67 BPU.scala 188:14]
  wire [2:0] _GEN_365 = _T_16 ? _GEN_316 : 3'h0; // @[Conditional.scala 39:67 BPU.scala 190:18]
  wire [24:0] _GEN_366 = _T_16 ? _GEN_317 : 25'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_367 = _T_16 ? _GEN_318 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_368 = _T_16 ? _GEN_319 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [31:0] _GEN_369 = _T_16 ? _GEN_320 : 32'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire  _GEN_370 = _T_16 & _GEN_321; // @[Conditional.scala 39:67 BPU.scala 188:14]
  wire [2:0] _GEN_371 = _T_16 ? _GEN_322 : 3'h0; // @[Conditional.scala 39:67 BPU.scala 190:18]
  wire [24:0] _GEN_372 = _T_16 ? _GEN_323 : 25'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_373 = _T_16 ? _GEN_324 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [1:0] _GEN_374 = _T_16 ? _GEN_325 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire [31:0] _GEN_375 = _T_16 ? _GEN_326 : 32'h0; // @[Conditional.scala 39:67 BPU.scala 191:13]
  wire  _GEN_376 = _T_16 & _T_23; // @[Conditional.scala 39:67 BPU.scala 203:15]
  wire [31:0] _GEN_377 = _T_16 ? _GEN_329 : 32'h0; // @[Conditional.scala 39:67 BPU.scala 205:17]
  wire  _GEN_378 = _T_16 & _GEN_330; // @[Conditional.scala 39:67 BPU.scala 204:14]
  wire [2:0] _GEN_379 = _T_16 ? 3'h0 : _GEN_344; // @[Conditional.scala 39:67 BPU.scala 189:18]
  wire [2:0] _GEN_384 = _T_14 ? _GEN_265 : _GEN_379; // @[Conditional.scala 40:58]
  wire  _GEN_415 = _T_14 ? 1'h0 : _GEN_376; // @[Conditional.scala 40:58 BPU.scala 203:15]
  wire [31:0] _GEN_416 = _T_14 ? 32'h0 : _GEN_377; // @[Conditional.scala 40:58 BPU.scala 205:17]
  wire  _GEN_417 = _T_14 ? 1'h0 : _GEN_378; // @[Conditional.scala 40:58 BPU.scala 204:14]
  wire  _bp_static_target_T_1 = ~ifu_pc_reg[31]; // @[BPU.scala 158:35]
  wire [31:0] _bp_static_target_T_3 = ifu_pc_reg + 32'h4; // @[BPU.scala 353:67]
  wire [27:0] bp_static_target_hi = ifu_pc_reg[31:4]; // @[BPU.scala 353:88]
  wire [31:0] _bp_static_target_T_4 = {bp_static_target_hi,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _bp_static_target_T_6 = _bp_static_target_T_4 + 32'h10; // @[BPU.scala 353:111]
  wire [31:0] bp_static_target = _bp_static_target_T_1 ? _bp_static_target_T_3 : _bp_static_target_T_6; // @[BPU.scala 353:26]
  wire  _T_28 = 2'h0 == ifu_state; // @[Conditional.scala 37:30]
  wire  _T_29 = ~io_ifu_is_reflush; // @[BPU.scala 361:26]
  wire  _T_30 = io_ifu_valid & ~io_ifu_is_reflush; // @[BPU.scala 361:23]
  wire [2:0] _GEN_420 = io_ifu_valid & ~io_ifu_is_reflush ? io_ifu_pc[6:4] : _GEN_384; // @[BPU.scala 361:43 BPU.scala 364:29]
  wire  _T_31 = 2'h1 == ifu_state; // @[Conditional.scala 37:30]
  wire [1:0] offset_0 = btb_0_io_out_offset;
  wire [3:0] _GEN_615 = {offset_0, 2'h0}; // @[BPU.scala 378:39]
  wire [4:0] _offset_real_T = {{1'd0}, _GEN_615}; // @[BPU.scala 378:39]
  wire  _bp_taken_T_3 = ifu_pc_reg[3:2] == offset_0; // @[BPU.scala 380:42]
  wire  _bp_taken_T_5 = ifu_pc_reg[3:2] <= offset_0; // @[BPU.scala 381:42]
  wire  _bp_taken_T_6 = _bp_static_target_T_1 ? _bp_taken_T_3 : _bp_taken_T_5; // @[BPU.scala 379:32]
  wire [1:0] btb_type_0 = btb_0_io_out_btb_type;
  wire [31:0] target_0 = btb_0_io_out_target;
  wire [31:0] _io_ifu_bp_target_T = io_ifu_bp_taken ? target_0 : bp_static_target; // @[BPU.scala 385:38]
  wire [1:0] offset_3 = btb_3_io_out_offset;
  wire [3:0] _GEN_616 = {offset_3, 2'h0}; // @[BPU.scala 378:39]
  wire [4:0] _offset_real_T_3 = {{1'd0}, _GEN_616}; // @[BPU.scala 378:39]
  wire [1:0] offset_2 = btb_2_io_out_offset;
  wire [3:0] _GEN_617 = {offset_2, 2'h0}; // @[BPU.scala 378:39]
  wire [4:0] _offset_real_T_2 = {{1'd0}, _GEN_617}; // @[BPU.scala 378:39]
  wire [1:0] offset_1 = btb_1_io_out_offset;
  wire [3:0] _GEN_618 = {offset_1, 2'h0}; // @[BPU.scala 378:39]
  wire [4:0] _offset_real_T_1 = {{1'd0}, _GEN_618}; // @[BPU.scala 378:39]
  wire [4:0] _GEN_441 = ifu_hit_0 ? _offset_real_T : 5'h0; // @[BPU.scala 375:29 BPU.scala 378:25]
  wire [4:0] _GEN_466 = ifu_hit_1 ? _offset_real_T_1 : _GEN_441; // @[BPU.scala 375:29 BPU.scala 378:25]
  wire [4:0] _GEN_491 = ifu_hit_2 ? _offset_real_T_2 : _GEN_466; // @[BPU.scala 375:29 BPU.scala 378:25]
  wire [4:0] _GEN_516 = ifu_hit_3 ? _offset_real_T_3 : _GEN_491; // @[BPU.scala 375:29 BPU.scala 378:25]
  wire [4:0] _GEN_526 = ifu_btb_hit & _T_29 ? _GEN_516 : 5'h0; // @[BPU.scala 373:45]
  wire [4:0] _GEN_554 = _T_31 ? _GEN_526 : 5'h0; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_575 = _T_28 ? 5'h0 : _GEN_554; // @[Conditional.scala 40:58]
  wire [3:0] offset_real = _GEN_575[3:0];
  wire [31:0] _GEN_619 = {{28'd0}, offset_real}; // @[BPU.scala 387:70]
  wire [31:0] _ras_io_addr_w_T_4 = _bp_static_target_T_4 + _GEN_619; // @[BPU.scala 387:70]
  wire [31:0] _ras_io_addr_w_T_6 = _ras_io_addr_w_T_4 + 32'h4; // @[BPU.scala 387:85]
  wire [31:0] _io_ifu_bp_target_T_1 = io_ifu_bp_taken ? ras_io_addr_r : bp_static_target; // @[BPU.scala 391:38]
  wire  _bp_taken_T_27 = ifu_pc_reg[3:2] == offset_3; // @[BPU.scala 380:42]
  wire  _bp_taken_T_29 = ifu_pc_reg[3:2] <= offset_3; // @[BPU.scala 381:42]
  wire  _bp_taken_T_30 = _bp_static_target_T_1 ? _bp_taken_T_27 : _bp_taken_T_29; // @[BPU.scala 379:32]
  wire  _bp_taken_T_19 = ifu_pc_reg[3:2] == offset_2; // @[BPU.scala 380:42]
  wire  _bp_taken_T_21 = ifu_pc_reg[3:2] <= offset_2; // @[BPU.scala 381:42]
  wire  _bp_taken_T_22 = _bp_static_target_T_1 ? _bp_taken_T_19 : _bp_taken_T_21; // @[BPU.scala 379:32]
  wire  _bp_taken_T_11 = ifu_pc_reg[3:2] == offset_1; // @[BPU.scala 380:42]
  wire  _bp_taken_T_13 = ifu_pc_reg[3:2] <= offset_1; // @[BPU.scala 381:42]
  wire  _bp_taken_T_14 = _bp_static_target_T_1 ? _bp_taken_T_11 : _bp_taken_T_13; // @[BPU.scala 379:32]
  wire  _GEN_467 = ifu_hit_1 ? _bp_taken_T_14 : ifu_hit_0 & _bp_taken_T_6; // @[BPU.scala 375:29 BPU.scala 379:22]
  wire  _GEN_492 = ifu_hit_2 ? _bp_taken_T_22 : _GEN_467; // @[BPU.scala 375:29 BPU.scala 379:22]
  wire  _GEN_517 = ifu_hit_3 ? _bp_taken_T_30 : _GEN_492; // @[BPU.scala 375:29 BPU.scala 379:22]
  wire  _GEN_527 = ifu_btb_hit & _T_29 & _GEN_517; // @[BPU.scala 373:45]
  wire  _GEN_555 = _T_31 & _GEN_527; // @[Conditional.scala 39:67]
  wire  bp_taken = _T_28 ? 1'h0 : _GEN_555; // @[Conditional.scala 40:58]
  wire  _GEN_424 = btb_type_0 == 2'h3 & bp_taken; // @[BPU.scala 396:52 BPU.scala 397:31 BPU.scala 352:19]
  wire [31:0] _GEN_425 = btb_type_0 == 2'h3 ? _io_ifu_bp_target_T : bp_static_target; // @[BPU.scala 396:52 BPU.scala 398:32 BPU.scala 354:20]
  wire [3:0] _GEN_426 = btb_type_0 == 2'h2 ? ifu_pc_reg[7:4] : 4'h0; // @[BPU.scala 392:54 BPU.scala 393:30 BPU.scala 199:18]
  wire  _GEN_427 = btb_type_0 == 2'h2 ? bp_taken & pht_io_br_taken : _GEN_424; // @[BPU.scala 392:54 BPU.scala 394:31]
  wire [31:0] _GEN_428 = btb_type_0 == 2'h2 ? _io_ifu_bp_target_T : _GEN_425; // @[BPU.scala 392:54 BPU.scala 395:32]
  wire  _GEN_429 = btb_type_0 == 2'h1 ? bp_taken : _GEN_427; // @[BPU.scala 388:51 BPU.scala 389:31]
  wire  _GEN_430 = btb_type_0 == 2'h1 ? bp_taken : _GEN_417; // @[BPU.scala 388:51 BPU.scala 390:26]
  wire [31:0] _GEN_431 = btb_type_0 == 2'h1 ? _io_ifu_bp_target_T_1 : _GEN_428; // @[BPU.scala 388:51 BPU.scala 391:32]
  wire [3:0] _GEN_432 = btb_type_0 == 2'h1 ? 4'h0 : _GEN_426; // @[BPU.scala 388:51 BPU.scala 199:18]
  wire  _GEN_433 = btb_type_0 == 2'h0 ? bp_taken : _GEN_429; // @[BPU.scala 383:45 BPU.scala 384:31]
  wire [31:0] _GEN_434 = btb_type_0 == 2'h0 ? _io_ifu_bp_target_T : _GEN_431; // @[BPU.scala 383:45 BPU.scala 385:32]
  wire  _GEN_435 = btb_type_0 == 2'h0 ? bp_taken : _GEN_415; // @[BPU.scala 383:45 BPU.scala 386:27]
  wire [31:0] _GEN_436 = btb_type_0 == 2'h0 ? _ras_io_addr_w_T_6 : _GEN_416; // @[BPU.scala 383:45 BPU.scala 387:29]
  wire  _GEN_437 = btb_type_0 == 2'h0 ? _GEN_417 : _GEN_430; // @[BPU.scala 383:45]
  wire [3:0] _GEN_438 = btb_type_0 == 2'h0 ? 4'h0 : _GEN_432; // @[BPU.scala 383:45 BPU.scala 199:18]
  wire [1:0] _GEN_439 = ifu_hit_0 ? btb_type_0 : 2'h3; // @[BPU.scala 375:29 BPU.scala 376:28 BPU.scala 357:18]
  wire [1:0] _GEN_440 = ifu_hit_0 ? offset_0 : 2'h0; // @[BPU.scala 375:29 BPU.scala 377:30 BPU.scala 355:20]
  wire  _GEN_443 = ifu_hit_0 & _GEN_433; // @[BPU.scala 375:29 BPU.scala 352:19]
  wire [31:0] _GEN_444 = ifu_hit_0 ? _GEN_434 : bp_static_target; // @[BPU.scala 375:29 BPU.scala 354:20]
  wire  _GEN_445 = ifu_hit_0 ? _GEN_435 : _GEN_415; // @[BPU.scala 375:29]
  wire [31:0] _GEN_446 = ifu_hit_0 ? _GEN_436 : _GEN_416; // @[BPU.scala 375:29]
  wire  _GEN_447 = ifu_hit_0 ? _GEN_437 : _GEN_417; // @[BPU.scala 375:29]
  wire [3:0] _GEN_448 = ifu_hit_0 ? _GEN_438 : 4'h0; // @[BPU.scala 375:29 BPU.scala 199:18]
  wire [1:0] btb_type_1 = btb_1_io_out_btb_type;
  wire [31:0] target_1 = btb_1_io_out_target;
  wire [31:0] _io_ifu_bp_target_T_4 = io_ifu_bp_taken ? target_1 : bp_static_target; // @[BPU.scala 385:38]
  wire  _GEN_449 = btb_type_1 == 2'h3 ? bp_taken : _GEN_443; // @[BPU.scala 396:52 BPU.scala 397:31]
  wire [31:0] _GEN_450 = btb_type_1 == 2'h3 ? _io_ifu_bp_target_T_4 : _GEN_444; // @[BPU.scala 396:52 BPU.scala 398:32]
  wire [3:0] _GEN_451 = btb_type_1 == 2'h2 ? ifu_pc_reg[7:4] : _GEN_448; // @[BPU.scala 392:54 BPU.scala 393:30]
  wire  _GEN_452 = btb_type_1 == 2'h2 ? bp_taken & pht_io_br_taken : _GEN_449; // @[BPU.scala 392:54 BPU.scala 394:31]
  wire [31:0] _GEN_453 = btb_type_1 == 2'h2 ? _io_ifu_bp_target_T_4 : _GEN_450; // @[BPU.scala 392:54 BPU.scala 395:32]
  wire  _GEN_454 = btb_type_1 == 2'h1 ? bp_taken : _GEN_452; // @[BPU.scala 388:51 BPU.scala 389:31]
  wire  _GEN_455 = btb_type_1 == 2'h1 ? bp_taken : _GEN_447; // @[BPU.scala 388:51 BPU.scala 390:26]
  wire [31:0] _GEN_456 = btb_type_1 == 2'h1 ? _io_ifu_bp_target_T_1 : _GEN_453; // @[BPU.scala 388:51 BPU.scala 391:32]
  wire [3:0] _GEN_457 = btb_type_1 == 2'h1 ? _GEN_448 : _GEN_451; // @[BPU.scala 388:51]
  wire  _GEN_458 = btb_type_1 == 2'h0 ? bp_taken : _GEN_454; // @[BPU.scala 383:45 BPU.scala 384:31]
  wire [31:0] _GEN_459 = btb_type_1 == 2'h0 ? _io_ifu_bp_target_T_4 : _GEN_456; // @[BPU.scala 383:45 BPU.scala 385:32]
  wire  _GEN_460 = btb_type_1 == 2'h0 ? bp_taken : _GEN_445; // @[BPU.scala 383:45 BPU.scala 386:27]
  wire [31:0] _GEN_461 = btb_type_1 == 2'h0 ? _ras_io_addr_w_T_6 : _GEN_446; // @[BPU.scala 383:45 BPU.scala 387:29]
  wire  _GEN_462 = btb_type_1 == 2'h0 ? _GEN_447 : _GEN_455; // @[BPU.scala 383:45]
  wire [3:0] _GEN_463 = btb_type_1 == 2'h0 ? _GEN_448 : _GEN_457; // @[BPU.scala 383:45]
  wire [1:0] _GEN_464 = ifu_hit_1 ? btb_type_1 : _GEN_439; // @[BPU.scala 375:29 BPU.scala 376:28]
  wire [1:0] _GEN_465 = ifu_hit_1 ? offset_1 : _GEN_440; // @[BPU.scala 375:29 BPU.scala 377:30]
  wire  _GEN_468 = ifu_hit_1 ? _GEN_458 : _GEN_443; // @[BPU.scala 375:29]
  wire [31:0] _GEN_469 = ifu_hit_1 ? _GEN_459 : _GEN_444; // @[BPU.scala 375:29]
  wire  _GEN_470 = ifu_hit_1 ? _GEN_460 : _GEN_445; // @[BPU.scala 375:29]
  wire [31:0] _GEN_471 = ifu_hit_1 ? _GEN_461 : _GEN_446; // @[BPU.scala 375:29]
  wire  _GEN_472 = ifu_hit_1 ? _GEN_462 : _GEN_447; // @[BPU.scala 375:29]
  wire [3:0] _GEN_473 = ifu_hit_1 ? _GEN_463 : _GEN_448; // @[BPU.scala 375:29]
  wire [1:0] btb_type_2 = btb_2_io_out_btb_type;
  wire [31:0] target_2 = btb_2_io_out_target;
  wire [31:0] _io_ifu_bp_target_T_8 = io_ifu_bp_taken ? target_2 : bp_static_target; // @[BPU.scala 385:38]
  wire  _GEN_474 = btb_type_2 == 2'h3 ? bp_taken : _GEN_468; // @[BPU.scala 396:52 BPU.scala 397:31]
  wire [31:0] _GEN_475 = btb_type_2 == 2'h3 ? _io_ifu_bp_target_T_8 : _GEN_469; // @[BPU.scala 396:52 BPU.scala 398:32]
  wire [3:0] _GEN_476 = btb_type_2 == 2'h2 ? ifu_pc_reg[7:4] : _GEN_473; // @[BPU.scala 392:54 BPU.scala 393:30]
  wire  _GEN_477 = btb_type_2 == 2'h2 ? bp_taken & pht_io_br_taken : _GEN_474; // @[BPU.scala 392:54 BPU.scala 394:31]
  wire [31:0] _GEN_478 = btb_type_2 == 2'h2 ? _io_ifu_bp_target_T_8 : _GEN_475; // @[BPU.scala 392:54 BPU.scala 395:32]
  wire  _GEN_479 = btb_type_2 == 2'h1 ? bp_taken : _GEN_477; // @[BPU.scala 388:51 BPU.scala 389:31]
  wire  _GEN_480 = btb_type_2 == 2'h1 ? bp_taken : _GEN_472; // @[BPU.scala 388:51 BPU.scala 390:26]
  wire [31:0] _GEN_481 = btb_type_2 == 2'h1 ? _io_ifu_bp_target_T_1 : _GEN_478; // @[BPU.scala 388:51 BPU.scala 391:32]
  wire [3:0] _GEN_482 = btb_type_2 == 2'h1 ? _GEN_473 : _GEN_476; // @[BPU.scala 388:51]
  wire  _GEN_483 = btb_type_2 == 2'h0 ? bp_taken : _GEN_479; // @[BPU.scala 383:45 BPU.scala 384:31]
  wire [31:0] _GEN_484 = btb_type_2 == 2'h0 ? _io_ifu_bp_target_T_8 : _GEN_481; // @[BPU.scala 383:45 BPU.scala 385:32]
  wire  _GEN_485 = btb_type_2 == 2'h0 ? bp_taken : _GEN_470; // @[BPU.scala 383:45 BPU.scala 386:27]
  wire [31:0] _GEN_486 = btb_type_2 == 2'h0 ? _ras_io_addr_w_T_6 : _GEN_471; // @[BPU.scala 383:45 BPU.scala 387:29]
  wire  _GEN_487 = btb_type_2 == 2'h0 ? _GEN_472 : _GEN_480; // @[BPU.scala 383:45]
  wire [3:0] _GEN_488 = btb_type_2 == 2'h0 ? _GEN_473 : _GEN_482; // @[BPU.scala 383:45]
  wire [1:0] _GEN_489 = ifu_hit_2 ? btb_type_2 : _GEN_464; // @[BPU.scala 375:29 BPU.scala 376:28]
  wire [1:0] _GEN_490 = ifu_hit_2 ? offset_2 : _GEN_465; // @[BPU.scala 375:29 BPU.scala 377:30]
  wire  _GEN_493 = ifu_hit_2 ? _GEN_483 : _GEN_468; // @[BPU.scala 375:29]
  wire [31:0] _GEN_494 = ifu_hit_2 ? _GEN_484 : _GEN_469; // @[BPU.scala 375:29]
  wire  _GEN_495 = ifu_hit_2 ? _GEN_485 : _GEN_470; // @[BPU.scala 375:29]
  wire [31:0] _GEN_496 = ifu_hit_2 ? _GEN_486 : _GEN_471; // @[BPU.scala 375:29]
  wire  _GEN_497 = ifu_hit_2 ? _GEN_487 : _GEN_472; // @[BPU.scala 375:29]
  wire [3:0] _GEN_498 = ifu_hit_2 ? _GEN_488 : _GEN_473; // @[BPU.scala 375:29]
  wire [1:0] btb_type_3 = btb_3_io_out_btb_type;
  wire [31:0] target_3 = btb_3_io_out_target;
  wire [31:0] _io_ifu_bp_target_T_12 = io_ifu_bp_taken ? target_3 : bp_static_target; // @[BPU.scala 385:38]
  wire  _GEN_499 = btb_type_3 == 2'h3 ? bp_taken : _GEN_493; // @[BPU.scala 396:52 BPU.scala 397:31]
  wire [31:0] _GEN_500 = btb_type_3 == 2'h3 ? _io_ifu_bp_target_T_12 : _GEN_494; // @[BPU.scala 396:52 BPU.scala 398:32]
  wire [3:0] _GEN_501 = btb_type_3 == 2'h2 ? ifu_pc_reg[7:4] : _GEN_498; // @[BPU.scala 392:54 BPU.scala 393:30]
  wire  _GEN_502 = btb_type_3 == 2'h2 ? bp_taken & pht_io_br_taken : _GEN_499; // @[BPU.scala 392:54 BPU.scala 394:31]
  wire [31:0] _GEN_503 = btb_type_3 == 2'h2 ? _io_ifu_bp_target_T_12 : _GEN_500; // @[BPU.scala 392:54 BPU.scala 395:32]
  wire  _GEN_504 = btb_type_3 == 2'h1 ? bp_taken : _GEN_502; // @[BPU.scala 388:51 BPU.scala 389:31]
  wire  _GEN_505 = btb_type_3 == 2'h1 ? bp_taken : _GEN_497; // @[BPU.scala 388:51 BPU.scala 390:26]
  wire [31:0] _GEN_506 = btb_type_3 == 2'h1 ? _io_ifu_bp_target_T_1 : _GEN_503; // @[BPU.scala 388:51 BPU.scala 391:32]
  wire [3:0] _GEN_507 = btb_type_3 == 2'h1 ? _GEN_498 : _GEN_501; // @[BPU.scala 388:51]
  wire  _GEN_508 = btb_type_3 == 2'h0 ? bp_taken : _GEN_504; // @[BPU.scala 383:45 BPU.scala 384:31]
  wire [31:0] _GEN_509 = btb_type_3 == 2'h0 ? _io_ifu_bp_target_T_12 : _GEN_506; // @[BPU.scala 383:45 BPU.scala 385:32]
  wire  _GEN_510 = btb_type_3 == 2'h0 ? bp_taken : _GEN_495; // @[BPU.scala 383:45 BPU.scala 386:27]
  wire [31:0] _GEN_511 = btb_type_3 == 2'h0 ? _ras_io_addr_w_T_6 : _GEN_496; // @[BPU.scala 383:45 BPU.scala 387:29]
  wire  _GEN_512 = btb_type_3 == 2'h0 ? _GEN_497 : _GEN_505; // @[BPU.scala 383:45]
  wire [3:0] _GEN_513 = btb_type_3 == 2'h0 ? _GEN_498 : _GEN_507; // @[BPU.scala 383:45]
  wire [1:0] _GEN_514 = ifu_hit_3 ? btb_type_3 : _GEN_489; // @[BPU.scala 375:29 BPU.scala 376:28]
  wire [1:0] _GEN_515 = ifu_hit_3 ? offset_3 : _GEN_490; // @[BPU.scala 375:29 BPU.scala 377:30]
  wire  _GEN_518 = ifu_hit_3 ? _GEN_508 : _GEN_493; // @[BPU.scala 375:29]
  wire [31:0] _GEN_519 = ifu_hit_3 ? _GEN_509 : _GEN_494; // @[BPU.scala 375:29]
  wire  _GEN_520 = ifu_hit_3 ? _GEN_510 : _GEN_495; // @[BPU.scala 375:29]
  wire [31:0] _GEN_521 = ifu_hit_3 ? _GEN_511 : _GEN_496; // @[BPU.scala 375:29]
  wire  _GEN_522 = ifu_hit_3 ? _GEN_512 : _GEN_497; // @[BPU.scala 375:29]
  wire [3:0] _GEN_523 = ifu_hit_3 ? _GEN_513 : _GEN_498; // @[BPU.scala 375:29]
  wire [1:0] _GEN_524 = ifu_btb_hit & _T_29 ? _GEN_514 : 2'h3; // @[BPU.scala 373:45 BPU.scala 357:18]
  wire [1:0] _GEN_525 = ifu_btb_hit & _T_29 ? _GEN_515 : 2'h0; // @[BPU.scala 373:45 BPU.scala 355:20]
  wire  _GEN_528 = ifu_btb_hit & _T_29 & _GEN_518; // @[BPU.scala 373:45 BPU.scala 403:25]
  wire [31:0] _GEN_529 = ifu_btb_hit & _T_29 ? _GEN_519 : bp_static_target; // @[BPU.scala 373:45 BPU.scala 404:26]
  wire  _GEN_530 = ifu_btb_hit & _T_29 ? _GEN_520 : _GEN_415; // @[BPU.scala 373:45]
  wire [31:0] _GEN_531 = ifu_btb_hit & _T_29 ? _GEN_521 : _GEN_416; // @[BPU.scala 373:45]
  wire  _GEN_532 = ifu_btb_hit & _T_29 ? _GEN_522 : _GEN_417; // @[BPU.scala 373:45]
  wire [3:0] _GEN_533 = ifu_btb_hit & _T_29 ? _GEN_523 : 4'h0; // @[BPU.scala 373:45 BPU.scala 199:18]
  wire [1:0] _GEN_534 = io_ifu_valid ? 2'h2 : 2'h0; // @[BPU.scala 412:31 BPU.scala 413:19 BPU.scala 415:19]
  wire [1:0] _GEN_535 = _T_30 ? 2'h1 : _GEN_534; // @[BPU.scala 407:43 BPU.scala 408:19]
  wire  _T_52 = 2'h2 == ifu_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_547 = _T_52 ? _GEN_420 : _GEN_384; // @[Conditional.scala 39:67]
  wire  _GEN_551 = _T_31 | _T_52; // @[Conditional.scala 39:67 BPU.scala 371:20]
  wire [1:0] _GEN_552 = _T_31 ? _GEN_524 : 2'h3; // @[Conditional.scala 39:67 BPU.scala 357:18]
  wire [1:0] _GEN_553 = _T_31 ? _GEN_525 : 2'h0; // @[Conditional.scala 39:67 BPU.scala 355:20]
  wire  _GEN_556 = _T_31 & _GEN_528; // @[Conditional.scala 39:67 BPU.scala 352:19]
  wire [31:0] _GEN_557 = _T_31 ? _GEN_529 : bp_static_target; // @[Conditional.scala 39:67 BPU.scala 354:20]
  wire  _GEN_558 = _T_31 ? _GEN_530 : _GEN_415; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_559 = _T_31 ? _GEN_531 : _GEN_416; // @[Conditional.scala 39:67]
  wire  _GEN_560 = _T_31 ? _GEN_532 : _GEN_417; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_561 = _T_31 ? _GEN_533 : 4'h0; // @[Conditional.scala 39:67 BPU.scala 199:18]
  wire [2:0] _GEN_563 = _T_31 ? _GEN_420 : _GEN_547; // @[Conditional.scala 39:67]
  BTB btb_0 ( // @[BPU.scala 183:21]
    .clock(btb_0_clock),
    .reset(btb_0_reset),
    .io_wen(btb_0_io_wen),
    .io_index_r(btb_0_io_index_r),
    .io_index_w(btb_0_io_index_w),
    .io_in_tag(btb_0_io_in_tag),
    .io_in_offset(btb_0_io_in_offset),
    .io_in_btb_type(btb_0_io_in_btb_type),
    .io_in_target(btb_0_io_in_target),
    .io_out_tag(btb_0_io_out_tag),
    .io_out_offset(btb_0_io_out_offset),
    .io_out_btb_type(btb_0_io_out_btb_type),
    .io_out_target(btb_0_io_out_target),
    .io_valid_r(btb_0_io_valid_r),
    .io_fence(btb_0_io_fence)
  );
  BTB btb_1 ( // @[BPU.scala 183:21]
    .clock(btb_1_clock),
    .reset(btb_1_reset),
    .io_wen(btb_1_io_wen),
    .io_index_r(btb_1_io_index_r),
    .io_index_w(btb_1_io_index_w),
    .io_in_tag(btb_1_io_in_tag),
    .io_in_offset(btb_1_io_in_offset),
    .io_in_btb_type(btb_1_io_in_btb_type),
    .io_in_target(btb_1_io_in_target),
    .io_out_tag(btb_1_io_out_tag),
    .io_out_offset(btb_1_io_out_offset),
    .io_out_btb_type(btb_1_io_out_btb_type),
    .io_out_target(btb_1_io_out_target),
    .io_valid_r(btb_1_io_valid_r),
    .io_fence(btb_1_io_fence)
  );
  BTB btb_2 ( // @[BPU.scala 183:21]
    .clock(btb_2_clock),
    .reset(btb_2_reset),
    .io_wen(btb_2_io_wen),
    .io_index_r(btb_2_io_index_r),
    .io_index_w(btb_2_io_index_w),
    .io_in_tag(btb_2_io_in_tag),
    .io_in_offset(btb_2_io_in_offset),
    .io_in_btb_type(btb_2_io_in_btb_type),
    .io_in_target(btb_2_io_in_target),
    .io_out_tag(btb_2_io_out_tag),
    .io_out_offset(btb_2_io_out_offset),
    .io_out_btb_type(btb_2_io_out_btb_type),
    .io_out_target(btb_2_io_out_target),
    .io_valid_r(btb_2_io_valid_r),
    .io_fence(btb_2_io_fence)
  );
  BTB btb_3 ( // @[BPU.scala 183:21]
    .clock(btb_3_clock),
    .reset(btb_3_reset),
    .io_wen(btb_3_io_wen),
    .io_index_r(btb_3_io_index_r),
    .io_index_w(btb_3_io_index_w),
    .io_in_tag(btb_3_io_in_tag),
    .io_in_offset(btb_3_io_in_offset),
    .io_in_btb_type(btb_3_io_in_btb_type),
    .io_in_target(btb_3_io_in_target),
    .io_out_tag(btb_3_io_out_tag),
    .io_out_offset(btb_3_io_out_offset),
    .io_out_btb_type(btb_3_io_out_btb_type),
    .io_out_target(btb_3_io_out_target),
    .io_valid_r(btb_3_io_valid_r),
    .io_fence(btb_3_io_fence)
  );
  PHT pht ( // @[BPU.scala 195:19]
    .clock(pht_clock),
    .reset(pht_reset),
    .io_inc(pht_io_inc),
    .io_dec(pht_io_dec),
    .io_index_w(pht_io_index_w),
    .io_index_r(pht_io_index_r),
    .io_fence(pht_io_fence),
    .io_br_taken(pht_io_br_taken)
  );
  RAS ras ( // @[BPU.scala 202:19]
    .clock(ras_clock),
    .reset(ras_reset),
    .io_call(ras_io_call),
    .io_ret(ras_io_ret),
    .io_call_count(ras_io_call_count),
    .io_ret_count(ras_io_ret_count),
    .io_addr_w(ras_io_addr_w),
    .io_addr_r(ras_io_addr_r),
    .io_reflush(ras_io_reflush),
    .io_fence(ras_io_fence)
  );
  assign io_ifu_bp_ok = _T_28 ? 1'h0 : _GEN_551; // @[Conditional.scala 40:58 BPU.scala 356:16]
  assign io_ifu_bp_taken = _T_28 ? 1'h0 : _GEN_556; // @[Conditional.scala 40:58 BPU.scala 352:19]
  assign io_ifu_bp_target = _T_28 ? bp_static_target : _GEN_557; // @[Conditional.scala 40:58 BPU.scala 354:20]
  assign io_ifu_bp_offset = _T_28 ? 2'h0 : _GEN_553; // @[Conditional.scala 40:58 BPU.scala 355:20]
  assign io_ifu_bp_type = _T_28 ? 2'h3 : _GEN_552; // @[Conditional.scala 40:58 BPU.scala 357:18]
  assign btb_0_clock = clock;
  assign btb_0_reset = reset;
  assign btb_0_io_wen = _T_14 ? 1'h0 : _GEN_352; // @[Conditional.scala 40:58 BPU.scala 188:14]
  assign btb_0_io_index_r = _T_28 ? _GEN_420 : _GEN_563; // @[Conditional.scala 40:58]
  assign btb_0_io_index_w = _T_14 ? 3'h0 : _GEN_353; // @[Conditional.scala 40:58 BPU.scala 190:18]
  assign btb_0_io_in_tag = _T_14 ? 25'h0 : _GEN_354; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_0_io_in_offset = _T_14 ? 2'h0 : _GEN_355; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_0_io_in_btb_type = _T_14 ? 2'h0 : _GEN_356; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_0_io_in_target = _T_14 ? 32'h0 : _GEN_357; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_0_io_fence = io_exu_fence; // @[BPU.scala 192:16]
  assign btb_1_clock = clock;
  assign btb_1_reset = reset;
  assign btb_1_io_wen = _T_14 ? 1'h0 : _GEN_358; // @[Conditional.scala 40:58 BPU.scala 188:14]
  assign btb_1_io_index_r = _T_28 ? _GEN_420 : _GEN_563; // @[Conditional.scala 40:58]
  assign btb_1_io_index_w = _T_14 ? 3'h0 : _GEN_359; // @[Conditional.scala 40:58 BPU.scala 190:18]
  assign btb_1_io_in_tag = _T_14 ? 25'h0 : _GEN_360; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_1_io_in_offset = _T_14 ? 2'h0 : _GEN_361; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_1_io_in_btb_type = _T_14 ? 2'h0 : _GEN_362; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_1_io_in_target = _T_14 ? 32'h0 : _GEN_363; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_1_io_fence = io_exu_fence; // @[BPU.scala 192:16]
  assign btb_2_clock = clock;
  assign btb_2_reset = reset;
  assign btb_2_io_wen = _T_14 ? 1'h0 : _GEN_364; // @[Conditional.scala 40:58 BPU.scala 188:14]
  assign btb_2_io_index_r = _T_28 ? _GEN_420 : _GEN_563; // @[Conditional.scala 40:58]
  assign btb_2_io_index_w = _T_14 ? 3'h0 : _GEN_365; // @[Conditional.scala 40:58 BPU.scala 190:18]
  assign btb_2_io_in_tag = _T_14 ? 25'h0 : _GEN_366; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_2_io_in_offset = _T_14 ? 2'h0 : _GEN_367; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_2_io_in_btb_type = _T_14 ? 2'h0 : _GEN_368; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_2_io_in_target = _T_14 ? 32'h0 : _GEN_369; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_2_io_fence = io_exu_fence; // @[BPU.scala 192:16]
  assign btb_3_clock = clock;
  assign btb_3_reset = reset;
  assign btb_3_io_wen = _T_14 ? 1'h0 : _GEN_370; // @[Conditional.scala 40:58 BPU.scala 188:14]
  assign btb_3_io_index_r = _T_28 ? _GEN_420 : _GEN_563; // @[Conditional.scala 40:58]
  assign btb_3_io_index_w = _T_14 ? 3'h0 : _GEN_371; // @[Conditional.scala 40:58 BPU.scala 190:18]
  assign btb_3_io_in_tag = _T_14 ? 25'h0 : _GEN_372; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_3_io_in_offset = _T_14 ? 2'h0 : _GEN_373; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_3_io_in_btb_type = _T_14 ? 2'h0 : _GEN_374; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_3_io_in_target = _T_14 ? 32'h0 : _GEN_375; // @[Conditional.scala 40:58 BPU.scala 191:13]
  assign btb_3_io_fence = io_exu_fence; // @[BPU.scala 192:16]
  assign pht_clock = clock;
  assign pht_reset = reset;
  assign pht_io_inc = _T_14 ? 1'h0 : _GEN_349; // @[Conditional.scala 40:58 BPU.scala 196:14]
  assign pht_io_dec = _T_14 ? 1'h0 : _GEN_350; // @[Conditional.scala 40:58 BPU.scala 197:14]
  assign pht_io_index_w = _T_14 ? 4'h0 : _GEN_348; // @[Conditional.scala 40:58 BPU.scala 198:18]
  assign pht_io_index_r = _T_28 ? 4'h0 : _GEN_561; // @[Conditional.scala 40:58 BPU.scala 199:18]
  assign pht_io_fence = io_exu_fence; // @[BPU.scala 200:16]
  assign ras_clock = clock;
  assign ras_reset = reset;
  assign ras_io_call = _T_28 ? _GEN_415 : _GEN_558; // @[Conditional.scala 40:58]
  assign ras_io_ret = _T_28 ? _GEN_417 : _GEN_560; // @[Conditional.scala 40:58]
  assign ras_io_call_count = io_ifu_call_count - io_exu_call_count; // @[BPU.scala 208:39]
  assign ras_io_ret_count = io_ifu_ret_count - io_exu_ret_count; // @[BPU.scala 209:37]
  assign ras_io_addr_w = _T_28 ? _GEN_416 : _GEN_559; // @[Conditional.scala 40:58]
  assign ras_io_reflush = io_ifu_is_reflush; // @[BPU.scala 207:18]
  assign ras_io_fence = io_exu_fence; // @[BPU.scala 206:16]
  always @(posedge clock) begin
    if (reset) begin // @[BPU.scala 161:27]
      ifu_pc_reg <= 32'h0; // @[BPU.scala 161:27]
    end else if (io_ifu_valid) begin // @[BPU.scala 169:20]
      ifu_pc_reg <= io_ifu_pc; // @[BPU.scala 170:16]
    end
    if (reset) begin // @[BPU.scala 162:27]
      exu_pc_reg <= 32'h0; // @[BPU.scala 162:27]
    end else if (io_exu_valid) begin // @[BPU.scala 173:20]
      exu_pc_reg <= io_exu_pc; // @[BPU.scala 174:16]
    end
    if (reset) begin // @[BPU.scala 163:33]
      exu_bp_taken_reg <= 1'h0; // @[BPU.scala 163:33]
    end else if (io_exu_valid) begin // @[BPU.scala 173:20]
      exu_bp_taken_reg <= io_exu_bp_taken; // @[BPU.scala 175:22]
    end
    if (reset) begin // @[BPU.scala 164:34]
      exu_bp_target_reg <= 32'h0; // @[BPU.scala 164:34]
    end else if (io_exu_valid) begin // @[BPU.scala 173:20]
      exu_bp_target_reg <= io_exu_bp_target; // @[BPU.scala 176:23]
    end
    if (reset) begin // @[BPU.scala 165:32]
      exu_bp_type_reg <= 2'h0; // @[BPU.scala 165:32]
    end else if (io_exu_valid) begin // @[BPU.scala 173:20]
      exu_bp_type_reg <= io_exu_bp_type; // @[BPU.scala 177:21]
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_0 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h0 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_0 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_0 <= _GEN_95;
      end
    end else begin
      plru0_0 <= _GEN_95;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_1 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h1 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_1 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_1 <= _GEN_96;
      end
    end else begin
      plru0_1 <= _GEN_96;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_2 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h2 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_2 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_2 <= _GEN_97;
      end
    end else begin
      plru0_2 <= _GEN_97;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_3 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h3 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_3 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_3 <= _GEN_98;
      end
    end else begin
      plru0_3 <= _GEN_98;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_4 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h4 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_4 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_4 <= _GEN_99;
      end
    end else begin
      plru0_4 <= _GEN_99;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_5 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h5 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_5 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_5 <= _GEN_100;
      end
    end else begin
      plru0_5 <= _GEN_100;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_6 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h6 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_6 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_6 <= _GEN_101;
      end
    end else begin
      plru0_6 <= _GEN_101;
    end
    if (reset) begin // @[BPU.scala 216:22]
      plru0_7 <= 1'h0; // @[BPU.scala 216:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (3'h7 == ifu_pc_reg[6:4]) begin // @[BPU.scala 261:38]
        plru0_7 <= ifu_hit_0 | ifu_hit_1; // @[BPU.scala 261:38]
      end else begin
        plru0_7 <= _GEN_102;
      end
    end else begin
      plru0_7 <= _GEN_102;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_0 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_0 <= _GEN_127;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_0 <= _GEN_135;
      end else begin
        plru1_0 <= _GEN_103;
      end
    end else begin
      plru1_0 <= _GEN_103;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_1 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_1 <= _GEN_128;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_1 <= _GEN_136;
      end else begin
        plru1_1 <= _GEN_104;
      end
    end else begin
      plru1_1 <= _GEN_104;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_2 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_2 <= _GEN_129;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_2 <= _GEN_137;
      end else begin
        plru1_2 <= _GEN_105;
      end
    end else begin
      plru1_2 <= _GEN_105;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_3 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_3 <= _GEN_130;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_3 <= _GEN_138;
      end else begin
        plru1_3 <= _GEN_106;
      end
    end else begin
      plru1_3 <= _GEN_106;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_4 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_4 <= _GEN_131;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_4 <= _GEN_139;
      end else begin
        plru1_4 <= _GEN_107;
      end
    end else begin
      plru1_4 <= _GEN_107;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_5 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_5 <= _GEN_132;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_5 <= _GEN_140;
      end else begin
        plru1_5 <= _GEN_108;
      end
    end else begin
      plru1_5 <= _GEN_108;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_6 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_6 <= _GEN_133;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_6 <= _GEN_141;
      end else begin
        plru1_6 <= _GEN_109;
      end
    end else begin
      plru1_6 <= _GEN_109;
    end
    if (reset) begin // @[BPU.scala 217:22]
      plru1_7 <= 1'h0; // @[BPU.scala 217:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru1_7 <= _GEN_134;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru1_7 <= _GEN_142;
      end else begin
        plru1_7 <= _GEN_110;
      end
    end else begin
      plru1_7 <= _GEN_110;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_0 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_0 <= _GEN_111;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_0 <= _GEN_111;
      end else begin
        plru2_0 <= _GEN_167;
      end
    end else begin
      plru2_0 <= _GEN_111;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_1 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_1 <= _GEN_112;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_1 <= _GEN_112;
      end else begin
        plru2_1 <= _GEN_168;
      end
    end else begin
      plru2_1 <= _GEN_112;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_2 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_2 <= _GEN_113;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_2 <= _GEN_113;
      end else begin
        plru2_2 <= _GEN_169;
      end
    end else begin
      plru2_2 <= _GEN_113;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_3 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_3 <= _GEN_114;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_3 <= _GEN_114;
      end else begin
        plru2_3 <= _GEN_170;
      end
    end else begin
      plru2_3 <= _GEN_114;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_4 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_4 <= _GEN_115;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_4 <= _GEN_115;
      end else begin
        plru2_4 <= _GEN_171;
      end
    end else begin
      plru2_4 <= _GEN_115;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_5 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_5 <= _GEN_116;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_5 <= _GEN_116;
      end else begin
        plru2_5 <= _GEN_172;
      end
    end else begin
      plru2_5 <= _GEN_116;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_6 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_6 <= _GEN_117;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_6 <= _GEN_117;
      end else begin
        plru2_6 <= _GEN_173;
      end
    end else begin
      plru2_6 <= _GEN_117;
    end
    if (reset) begin // @[BPU.scala 218:22]
      plru2_7 <= 1'h0; // @[BPU.scala 218:22]
    end else if (ifu_state == 2'h1 & ifu_btb_hit) begin // @[BPU.scala 260:52]
      if (ifu_hit_0) begin // @[BPU.scala 262:23]
        plru2_7 <= _GEN_118;
      end else if (ifu_hit_1) begin // @[BPU.scala 264:30]
        plru2_7 <= _GEN_118;
      end else begin
        plru2_7 <= _GEN_174;
      end
    end else begin
      plru2_7 <= _GEN_118;
    end
    if (reset) begin // @[BPU.scala 234:26]
      ifu_state <= 2'h0; // @[BPU.scala 234:26]
    end else if (_T_28) begin // @[Conditional.scala 40:58]
      if (io_ifu_valid & ~io_ifu_is_reflush) begin // @[BPU.scala 361:43]
        ifu_state <= 2'h1; // @[BPU.scala 362:19]
      end else if (io_ifu_valid) begin // @[BPU.scala 366:31]
        ifu_state <= 2'h2; // @[BPU.scala 367:19]
      end
    end else if (_T_31) begin // @[Conditional.scala 39:67]
      ifu_state <= _GEN_535;
    end else if (_T_52) begin // @[Conditional.scala 39:67]
      ifu_state <= _GEN_535;
    end
    if (reset) begin // @[BPU.scala 235:26]
      exu_state <= 2'h0; // @[BPU.scala 235:26]
    end else if (_T_14) begin // @[Conditional.scala 40:58]
      if (io_exu_valid & io_exu_bp_wrong) begin // @[BPU.scala 284:40]
        exu_state <= 2'h1; // @[BPU.scala 285:19]
      end else if (io_exu_valid) begin // @[BPU.scala 289:31]
        exu_state <= 2'h2; // @[BPU.scala 290:19]
      end
    end else if (_T_16) begin // @[Conditional.scala 39:67]
      exu_state <= 2'h0;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      exu_state <= _GEN_335;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ifu_pc_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  exu_pc_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  exu_bp_taken_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  exu_bp_target_reg = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  exu_bp_type_reg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  plru0_0 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  plru0_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  plru0_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  plru0_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  plru0_4 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  plru0_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  plru0_6 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  plru0_7 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  plru1_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  plru1_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  plru1_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  plru1_3 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  plru1_4 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  plru1_5 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  plru1_6 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  plru1_7 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  plru2_0 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  plru2_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  plru2_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  plru2_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  plru2_4 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  plru2_5 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  plru2_6 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  plru2_7 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  ifu_state = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  exu_state = _RAND_30[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module META(
  input         clock,
  input         reset,
  input  [5:0]  io_index,
  output [21:0] io_tag_r,
  input  [21:0] io_tag_w,
  input         io_tag_wen,
  output        io_dirty_r,
  input         io_dirty_w,
  input         io_dirty_wen,
  output        io_valid_r,
  input         io_fence,
  output        io_fence_dirty
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] tag [0:63]; // @[META.scala 20:24]
  wire [21:0] tag_io_tag_r_MPORT_data; // @[META.scala 20:24]
  wire [5:0] tag_io_tag_r_MPORT_addr; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_addr; // @[META.scala 20:24]
  wire  tag_MPORT_mask; // @[META.scala 20:24]
  wire  tag_MPORT_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_1_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_1_addr; // @[META.scala 20:24]
  wire  tag_MPORT_1_mask; // @[META.scala 20:24]
  wire  tag_MPORT_1_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_2_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_2_addr; // @[META.scala 20:24]
  wire  tag_MPORT_2_mask; // @[META.scala 20:24]
  wire  tag_MPORT_2_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_3_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_3_addr; // @[META.scala 20:24]
  wire  tag_MPORT_3_mask; // @[META.scala 20:24]
  wire  tag_MPORT_3_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_4_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_4_addr; // @[META.scala 20:24]
  wire  tag_MPORT_4_mask; // @[META.scala 20:24]
  wire  tag_MPORT_4_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_5_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_5_addr; // @[META.scala 20:24]
  wire  tag_MPORT_5_mask; // @[META.scala 20:24]
  wire  tag_MPORT_5_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_6_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_6_addr; // @[META.scala 20:24]
  wire  tag_MPORT_6_mask; // @[META.scala 20:24]
  wire  tag_MPORT_6_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_7_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_7_addr; // @[META.scala 20:24]
  wire  tag_MPORT_7_mask; // @[META.scala 20:24]
  wire  tag_MPORT_7_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_8_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_8_addr; // @[META.scala 20:24]
  wire  tag_MPORT_8_mask; // @[META.scala 20:24]
  wire  tag_MPORT_8_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_9_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_9_addr; // @[META.scala 20:24]
  wire  tag_MPORT_9_mask; // @[META.scala 20:24]
  wire  tag_MPORT_9_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_10_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_10_addr; // @[META.scala 20:24]
  wire  tag_MPORT_10_mask; // @[META.scala 20:24]
  wire  tag_MPORT_10_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_11_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_11_addr; // @[META.scala 20:24]
  wire  tag_MPORT_11_mask; // @[META.scala 20:24]
  wire  tag_MPORT_11_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_12_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_12_addr; // @[META.scala 20:24]
  wire  tag_MPORT_12_mask; // @[META.scala 20:24]
  wire  tag_MPORT_12_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_13_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_13_addr; // @[META.scala 20:24]
  wire  tag_MPORT_13_mask; // @[META.scala 20:24]
  wire  tag_MPORT_13_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_14_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_14_addr; // @[META.scala 20:24]
  wire  tag_MPORT_14_mask; // @[META.scala 20:24]
  wire  tag_MPORT_14_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_15_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_15_addr; // @[META.scala 20:24]
  wire  tag_MPORT_15_mask; // @[META.scala 20:24]
  wire  tag_MPORT_15_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_16_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_16_addr; // @[META.scala 20:24]
  wire  tag_MPORT_16_mask; // @[META.scala 20:24]
  wire  tag_MPORT_16_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_17_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_17_addr; // @[META.scala 20:24]
  wire  tag_MPORT_17_mask; // @[META.scala 20:24]
  wire  tag_MPORT_17_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_18_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_18_addr; // @[META.scala 20:24]
  wire  tag_MPORT_18_mask; // @[META.scala 20:24]
  wire  tag_MPORT_18_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_19_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_19_addr; // @[META.scala 20:24]
  wire  tag_MPORT_19_mask; // @[META.scala 20:24]
  wire  tag_MPORT_19_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_20_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_20_addr; // @[META.scala 20:24]
  wire  tag_MPORT_20_mask; // @[META.scala 20:24]
  wire  tag_MPORT_20_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_21_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_21_addr; // @[META.scala 20:24]
  wire  tag_MPORT_21_mask; // @[META.scala 20:24]
  wire  tag_MPORT_21_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_22_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_22_addr; // @[META.scala 20:24]
  wire  tag_MPORT_22_mask; // @[META.scala 20:24]
  wire  tag_MPORT_22_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_23_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_23_addr; // @[META.scala 20:24]
  wire  tag_MPORT_23_mask; // @[META.scala 20:24]
  wire  tag_MPORT_23_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_24_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_24_addr; // @[META.scala 20:24]
  wire  tag_MPORT_24_mask; // @[META.scala 20:24]
  wire  tag_MPORT_24_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_25_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_25_addr; // @[META.scala 20:24]
  wire  tag_MPORT_25_mask; // @[META.scala 20:24]
  wire  tag_MPORT_25_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_26_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_26_addr; // @[META.scala 20:24]
  wire  tag_MPORT_26_mask; // @[META.scala 20:24]
  wire  tag_MPORT_26_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_27_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_27_addr; // @[META.scala 20:24]
  wire  tag_MPORT_27_mask; // @[META.scala 20:24]
  wire  tag_MPORT_27_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_28_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_28_addr; // @[META.scala 20:24]
  wire  tag_MPORT_28_mask; // @[META.scala 20:24]
  wire  tag_MPORT_28_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_29_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_29_addr; // @[META.scala 20:24]
  wire  tag_MPORT_29_mask; // @[META.scala 20:24]
  wire  tag_MPORT_29_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_30_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_30_addr; // @[META.scala 20:24]
  wire  tag_MPORT_30_mask; // @[META.scala 20:24]
  wire  tag_MPORT_30_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_31_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_31_addr; // @[META.scala 20:24]
  wire  tag_MPORT_31_mask; // @[META.scala 20:24]
  wire  tag_MPORT_31_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_32_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_32_addr; // @[META.scala 20:24]
  wire  tag_MPORT_32_mask; // @[META.scala 20:24]
  wire  tag_MPORT_32_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_33_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_33_addr; // @[META.scala 20:24]
  wire  tag_MPORT_33_mask; // @[META.scala 20:24]
  wire  tag_MPORT_33_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_34_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_34_addr; // @[META.scala 20:24]
  wire  tag_MPORT_34_mask; // @[META.scala 20:24]
  wire  tag_MPORT_34_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_35_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_35_addr; // @[META.scala 20:24]
  wire  tag_MPORT_35_mask; // @[META.scala 20:24]
  wire  tag_MPORT_35_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_36_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_36_addr; // @[META.scala 20:24]
  wire  tag_MPORT_36_mask; // @[META.scala 20:24]
  wire  tag_MPORT_36_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_37_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_37_addr; // @[META.scala 20:24]
  wire  tag_MPORT_37_mask; // @[META.scala 20:24]
  wire  tag_MPORT_37_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_38_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_38_addr; // @[META.scala 20:24]
  wire  tag_MPORT_38_mask; // @[META.scala 20:24]
  wire  tag_MPORT_38_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_39_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_39_addr; // @[META.scala 20:24]
  wire  tag_MPORT_39_mask; // @[META.scala 20:24]
  wire  tag_MPORT_39_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_40_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_40_addr; // @[META.scala 20:24]
  wire  tag_MPORT_40_mask; // @[META.scala 20:24]
  wire  tag_MPORT_40_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_41_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_41_addr; // @[META.scala 20:24]
  wire  tag_MPORT_41_mask; // @[META.scala 20:24]
  wire  tag_MPORT_41_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_42_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_42_addr; // @[META.scala 20:24]
  wire  tag_MPORT_42_mask; // @[META.scala 20:24]
  wire  tag_MPORT_42_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_43_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_43_addr; // @[META.scala 20:24]
  wire  tag_MPORT_43_mask; // @[META.scala 20:24]
  wire  tag_MPORT_43_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_44_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_44_addr; // @[META.scala 20:24]
  wire  tag_MPORT_44_mask; // @[META.scala 20:24]
  wire  tag_MPORT_44_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_45_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_45_addr; // @[META.scala 20:24]
  wire  tag_MPORT_45_mask; // @[META.scala 20:24]
  wire  tag_MPORT_45_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_46_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_46_addr; // @[META.scala 20:24]
  wire  tag_MPORT_46_mask; // @[META.scala 20:24]
  wire  tag_MPORT_46_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_47_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_47_addr; // @[META.scala 20:24]
  wire  tag_MPORT_47_mask; // @[META.scala 20:24]
  wire  tag_MPORT_47_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_48_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_48_addr; // @[META.scala 20:24]
  wire  tag_MPORT_48_mask; // @[META.scala 20:24]
  wire  tag_MPORT_48_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_49_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_49_addr; // @[META.scala 20:24]
  wire  tag_MPORT_49_mask; // @[META.scala 20:24]
  wire  tag_MPORT_49_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_50_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_50_addr; // @[META.scala 20:24]
  wire  tag_MPORT_50_mask; // @[META.scala 20:24]
  wire  tag_MPORT_50_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_51_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_51_addr; // @[META.scala 20:24]
  wire  tag_MPORT_51_mask; // @[META.scala 20:24]
  wire  tag_MPORT_51_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_52_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_52_addr; // @[META.scala 20:24]
  wire  tag_MPORT_52_mask; // @[META.scala 20:24]
  wire  tag_MPORT_52_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_53_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_53_addr; // @[META.scala 20:24]
  wire  tag_MPORT_53_mask; // @[META.scala 20:24]
  wire  tag_MPORT_53_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_54_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_54_addr; // @[META.scala 20:24]
  wire  tag_MPORT_54_mask; // @[META.scala 20:24]
  wire  tag_MPORT_54_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_55_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_55_addr; // @[META.scala 20:24]
  wire  tag_MPORT_55_mask; // @[META.scala 20:24]
  wire  tag_MPORT_55_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_56_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_56_addr; // @[META.scala 20:24]
  wire  tag_MPORT_56_mask; // @[META.scala 20:24]
  wire  tag_MPORT_56_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_57_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_57_addr; // @[META.scala 20:24]
  wire  tag_MPORT_57_mask; // @[META.scala 20:24]
  wire  tag_MPORT_57_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_58_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_58_addr; // @[META.scala 20:24]
  wire  tag_MPORT_58_mask; // @[META.scala 20:24]
  wire  tag_MPORT_58_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_59_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_59_addr; // @[META.scala 20:24]
  wire  tag_MPORT_59_mask; // @[META.scala 20:24]
  wire  tag_MPORT_59_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_60_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_60_addr; // @[META.scala 20:24]
  wire  tag_MPORT_60_mask; // @[META.scala 20:24]
  wire  tag_MPORT_60_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_61_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_61_addr; // @[META.scala 20:24]
  wire  tag_MPORT_61_mask; // @[META.scala 20:24]
  wire  tag_MPORT_61_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_62_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_62_addr; // @[META.scala 20:24]
  wire  tag_MPORT_62_mask; // @[META.scala 20:24]
  wire  tag_MPORT_62_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_63_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_63_addr; // @[META.scala 20:24]
  wire  tag_MPORT_63_mask; // @[META.scala 20:24]
  wire  tag_MPORT_63_en; // @[META.scala 20:24]
  wire [21:0] tag_MPORT_64_data; // @[META.scala 20:24]
  wire [5:0] tag_MPORT_64_addr; // @[META.scala 20:24]
  wire  tag_MPORT_64_mask; // @[META.scala 20:24]
  wire  tag_MPORT_64_en; // @[META.scala 20:24]
  reg [5:0] tag_io_tag_r_MPORT_addr_pipe_0;
  reg  valid_0; // @[META.scala 22:22]
  reg  valid_1; // @[META.scala 22:22]
  reg  valid_2; // @[META.scala 22:22]
  reg  valid_3; // @[META.scala 22:22]
  reg  valid_4; // @[META.scala 22:22]
  reg  valid_5; // @[META.scala 22:22]
  reg  valid_6; // @[META.scala 22:22]
  reg  valid_7; // @[META.scala 22:22]
  reg  valid_8; // @[META.scala 22:22]
  reg  valid_9; // @[META.scala 22:22]
  reg  valid_10; // @[META.scala 22:22]
  reg  valid_11; // @[META.scala 22:22]
  reg  valid_12; // @[META.scala 22:22]
  reg  valid_13; // @[META.scala 22:22]
  reg  valid_14; // @[META.scala 22:22]
  reg  valid_15; // @[META.scala 22:22]
  reg  valid_16; // @[META.scala 22:22]
  reg  valid_17; // @[META.scala 22:22]
  reg  valid_18; // @[META.scala 22:22]
  reg  valid_19; // @[META.scala 22:22]
  reg  valid_20; // @[META.scala 22:22]
  reg  valid_21; // @[META.scala 22:22]
  reg  valid_22; // @[META.scala 22:22]
  reg  valid_23; // @[META.scala 22:22]
  reg  valid_24; // @[META.scala 22:22]
  reg  valid_25; // @[META.scala 22:22]
  reg  valid_26; // @[META.scala 22:22]
  reg  valid_27; // @[META.scala 22:22]
  reg  valid_28; // @[META.scala 22:22]
  reg  valid_29; // @[META.scala 22:22]
  reg  valid_30; // @[META.scala 22:22]
  reg  valid_31; // @[META.scala 22:22]
  reg  valid_32; // @[META.scala 22:22]
  reg  valid_33; // @[META.scala 22:22]
  reg  valid_34; // @[META.scala 22:22]
  reg  valid_35; // @[META.scala 22:22]
  reg  valid_36; // @[META.scala 22:22]
  reg  valid_37; // @[META.scala 22:22]
  reg  valid_38; // @[META.scala 22:22]
  reg  valid_39; // @[META.scala 22:22]
  reg  valid_40; // @[META.scala 22:22]
  reg  valid_41; // @[META.scala 22:22]
  reg  valid_42; // @[META.scala 22:22]
  reg  valid_43; // @[META.scala 22:22]
  reg  valid_44; // @[META.scala 22:22]
  reg  valid_45; // @[META.scala 22:22]
  reg  valid_46; // @[META.scala 22:22]
  reg  valid_47; // @[META.scala 22:22]
  reg  valid_48; // @[META.scala 22:22]
  reg  valid_49; // @[META.scala 22:22]
  reg  valid_50; // @[META.scala 22:22]
  reg  valid_51; // @[META.scala 22:22]
  reg  valid_52; // @[META.scala 22:22]
  reg  valid_53; // @[META.scala 22:22]
  reg  valid_54; // @[META.scala 22:22]
  reg  valid_55; // @[META.scala 22:22]
  reg  valid_56; // @[META.scala 22:22]
  reg  valid_57; // @[META.scala 22:22]
  reg  valid_58; // @[META.scala 22:22]
  reg  valid_59; // @[META.scala 22:22]
  reg  valid_60; // @[META.scala 22:22]
  reg  valid_61; // @[META.scala 22:22]
  reg  valid_62; // @[META.scala 22:22]
  reg  valid_63; // @[META.scala 22:22]
  reg  dirty_0; // @[META.scala 23:22]
  reg  dirty_1; // @[META.scala 23:22]
  reg  dirty_2; // @[META.scala 23:22]
  reg  dirty_3; // @[META.scala 23:22]
  reg  dirty_4; // @[META.scala 23:22]
  reg  dirty_5; // @[META.scala 23:22]
  reg  dirty_6; // @[META.scala 23:22]
  reg  dirty_7; // @[META.scala 23:22]
  reg  dirty_8; // @[META.scala 23:22]
  reg  dirty_9; // @[META.scala 23:22]
  reg  dirty_10; // @[META.scala 23:22]
  reg  dirty_11; // @[META.scala 23:22]
  reg  dirty_12; // @[META.scala 23:22]
  reg  dirty_13; // @[META.scala 23:22]
  reg  dirty_14; // @[META.scala 23:22]
  reg  dirty_15; // @[META.scala 23:22]
  reg  dirty_16; // @[META.scala 23:22]
  reg  dirty_17; // @[META.scala 23:22]
  reg  dirty_18; // @[META.scala 23:22]
  reg  dirty_19; // @[META.scala 23:22]
  reg  dirty_20; // @[META.scala 23:22]
  reg  dirty_21; // @[META.scala 23:22]
  reg  dirty_22; // @[META.scala 23:22]
  reg  dirty_23; // @[META.scala 23:22]
  reg  dirty_24; // @[META.scala 23:22]
  reg  dirty_25; // @[META.scala 23:22]
  reg  dirty_26; // @[META.scala 23:22]
  reg  dirty_27; // @[META.scala 23:22]
  reg  dirty_28; // @[META.scala 23:22]
  reg  dirty_29; // @[META.scala 23:22]
  reg  dirty_30; // @[META.scala 23:22]
  reg  dirty_31; // @[META.scala 23:22]
  reg  dirty_32; // @[META.scala 23:22]
  reg  dirty_33; // @[META.scala 23:22]
  reg  dirty_34; // @[META.scala 23:22]
  reg  dirty_35; // @[META.scala 23:22]
  reg  dirty_36; // @[META.scala 23:22]
  reg  dirty_37; // @[META.scala 23:22]
  reg  dirty_38; // @[META.scala 23:22]
  reg  dirty_39; // @[META.scala 23:22]
  reg  dirty_40; // @[META.scala 23:22]
  reg  dirty_41; // @[META.scala 23:22]
  reg  dirty_42; // @[META.scala 23:22]
  reg  dirty_43; // @[META.scala 23:22]
  reg  dirty_44; // @[META.scala 23:22]
  reg  dirty_45; // @[META.scala 23:22]
  reg  dirty_46; // @[META.scala 23:22]
  reg  dirty_47; // @[META.scala 23:22]
  reg  dirty_48; // @[META.scala 23:22]
  reg  dirty_49; // @[META.scala 23:22]
  reg  dirty_50; // @[META.scala 23:22]
  reg  dirty_51; // @[META.scala 23:22]
  reg  dirty_52; // @[META.scala 23:22]
  reg  dirty_53; // @[META.scala 23:22]
  reg  dirty_54; // @[META.scala 23:22]
  reg  dirty_55; // @[META.scala 23:22]
  reg  dirty_56; // @[META.scala 23:22]
  reg  dirty_57; // @[META.scala 23:22]
  reg  dirty_58; // @[META.scala 23:22]
  reg  dirty_59; // @[META.scala 23:22]
  reg  dirty_60; // @[META.scala 23:22]
  reg  dirty_61; // @[META.scala 23:22]
  reg  dirty_62; // @[META.scala 23:22]
  reg  dirty_63; // @[META.scala 23:22]
  wire  _GEN_0 = 6'h0 == io_index | valid_0; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_1 = 6'h1 == io_index | valid_1; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_2 = 6'h2 == io_index | valid_2; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_3 = 6'h3 == io_index | valid_3; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_4 = 6'h4 == io_index | valid_4; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_5 = 6'h5 == io_index | valid_5; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_6 = 6'h6 == io_index | valid_6; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_7 = 6'h7 == io_index | valid_7; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_8 = 6'h8 == io_index | valid_8; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_9 = 6'h9 == io_index | valid_9; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_10 = 6'ha == io_index | valid_10; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_11 = 6'hb == io_index | valid_11; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_12 = 6'hc == io_index | valid_12; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_13 = 6'hd == io_index | valid_13; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_14 = 6'he == io_index | valid_14; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_15 = 6'hf == io_index | valid_15; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_16 = 6'h10 == io_index | valid_16; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_17 = 6'h11 == io_index | valid_17; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_18 = 6'h12 == io_index | valid_18; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_19 = 6'h13 == io_index | valid_19; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_20 = 6'h14 == io_index | valid_20; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_21 = 6'h15 == io_index | valid_21; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_22 = 6'h16 == io_index | valid_22; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_23 = 6'h17 == io_index | valid_23; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_24 = 6'h18 == io_index | valid_24; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_25 = 6'h19 == io_index | valid_25; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_26 = 6'h1a == io_index | valid_26; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_27 = 6'h1b == io_index | valid_27; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_28 = 6'h1c == io_index | valid_28; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_29 = 6'h1d == io_index | valid_29; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_30 = 6'h1e == io_index | valid_30; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_31 = 6'h1f == io_index | valid_31; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_32 = 6'h20 == io_index | valid_32; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_33 = 6'h21 == io_index | valid_33; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_34 = 6'h22 == io_index | valid_34; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_35 = 6'h23 == io_index | valid_35; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_36 = 6'h24 == io_index | valid_36; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_37 = 6'h25 == io_index | valid_37; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_38 = 6'h26 == io_index | valid_38; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_39 = 6'h27 == io_index | valid_39; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_40 = 6'h28 == io_index | valid_40; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_41 = 6'h29 == io_index | valid_41; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_42 = 6'h2a == io_index | valid_42; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_43 = 6'h2b == io_index | valid_43; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_44 = 6'h2c == io_index | valid_44; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_45 = 6'h2d == io_index | valid_45; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_46 = 6'h2e == io_index | valid_46; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_47 = 6'h2f == io_index | valid_47; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_48 = 6'h30 == io_index | valid_48; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_49 = 6'h31 == io_index | valid_49; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_50 = 6'h32 == io_index | valid_50; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_51 = 6'h33 == io_index | valid_51; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_52 = 6'h34 == io_index | valid_52; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_53 = 6'h35 == io_index | valid_53; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_54 = 6'h36 == io_index | valid_54; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_55 = 6'h37 == io_index | valid_55; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_56 = 6'h38 == io_index | valid_56; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_57 = 6'h39 == io_index | valid_57; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_58 = 6'h3a == io_index | valid_58; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_59 = 6'h3b == io_index | valid_59; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_60 = 6'h3c == io_index | valid_60; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_61 = 6'h3d == io_index | valid_61; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_62 = 6'h3e == io_index | valid_62; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  wire  _GEN_63 = 6'h3f == io_index | valid_63; // @[META.scala 27:18 META.scala 27:18 META.scala 22:22]
  reg  io_dirty_r_REG; // @[META.scala 31:24]
  wire  _GEN_134 = 6'h1 == io_index ? dirty_1 : dirty_0; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_135 = 6'h2 == io_index ? dirty_2 : _GEN_134; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_136 = 6'h3 == io_index ? dirty_3 : _GEN_135; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_137 = 6'h4 == io_index ? dirty_4 : _GEN_136; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_138 = 6'h5 == io_index ? dirty_5 : _GEN_137; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_139 = 6'h6 == io_index ? dirty_6 : _GEN_138; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_140 = 6'h7 == io_index ? dirty_7 : _GEN_139; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_141 = 6'h8 == io_index ? dirty_8 : _GEN_140; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_142 = 6'h9 == io_index ? dirty_9 : _GEN_141; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_143 = 6'ha == io_index ? dirty_10 : _GEN_142; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_144 = 6'hb == io_index ? dirty_11 : _GEN_143; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_145 = 6'hc == io_index ? dirty_12 : _GEN_144; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_146 = 6'hd == io_index ? dirty_13 : _GEN_145; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_147 = 6'he == io_index ? dirty_14 : _GEN_146; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_148 = 6'hf == io_index ? dirty_15 : _GEN_147; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_149 = 6'h10 == io_index ? dirty_16 : _GEN_148; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_150 = 6'h11 == io_index ? dirty_17 : _GEN_149; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_151 = 6'h12 == io_index ? dirty_18 : _GEN_150; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_152 = 6'h13 == io_index ? dirty_19 : _GEN_151; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_153 = 6'h14 == io_index ? dirty_20 : _GEN_152; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_154 = 6'h15 == io_index ? dirty_21 : _GEN_153; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_155 = 6'h16 == io_index ? dirty_22 : _GEN_154; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_156 = 6'h17 == io_index ? dirty_23 : _GEN_155; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_157 = 6'h18 == io_index ? dirty_24 : _GEN_156; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_158 = 6'h19 == io_index ? dirty_25 : _GEN_157; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_159 = 6'h1a == io_index ? dirty_26 : _GEN_158; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_160 = 6'h1b == io_index ? dirty_27 : _GEN_159; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_161 = 6'h1c == io_index ? dirty_28 : _GEN_160; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_162 = 6'h1d == io_index ? dirty_29 : _GEN_161; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_163 = 6'h1e == io_index ? dirty_30 : _GEN_162; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_164 = 6'h1f == io_index ? dirty_31 : _GEN_163; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_165 = 6'h20 == io_index ? dirty_32 : _GEN_164; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_166 = 6'h21 == io_index ? dirty_33 : _GEN_165; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_167 = 6'h22 == io_index ? dirty_34 : _GEN_166; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_168 = 6'h23 == io_index ? dirty_35 : _GEN_167; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_169 = 6'h24 == io_index ? dirty_36 : _GEN_168; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_170 = 6'h25 == io_index ? dirty_37 : _GEN_169; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_171 = 6'h26 == io_index ? dirty_38 : _GEN_170; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_172 = 6'h27 == io_index ? dirty_39 : _GEN_171; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_173 = 6'h28 == io_index ? dirty_40 : _GEN_172; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_174 = 6'h29 == io_index ? dirty_41 : _GEN_173; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_175 = 6'h2a == io_index ? dirty_42 : _GEN_174; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_176 = 6'h2b == io_index ? dirty_43 : _GEN_175; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_177 = 6'h2c == io_index ? dirty_44 : _GEN_176; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_178 = 6'h2d == io_index ? dirty_45 : _GEN_177; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_179 = 6'h2e == io_index ? dirty_46 : _GEN_178; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_180 = 6'h2f == io_index ? dirty_47 : _GEN_179; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_181 = 6'h30 == io_index ? dirty_48 : _GEN_180; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_182 = 6'h31 == io_index ? dirty_49 : _GEN_181; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_183 = 6'h32 == io_index ? dirty_50 : _GEN_182; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_184 = 6'h33 == io_index ? dirty_51 : _GEN_183; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_185 = 6'h34 == io_index ? dirty_52 : _GEN_184; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_186 = 6'h35 == io_index ? dirty_53 : _GEN_185; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_187 = 6'h36 == io_index ? dirty_54 : _GEN_186; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_188 = 6'h37 == io_index ? dirty_55 : _GEN_187; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_189 = 6'h38 == io_index ? dirty_56 : _GEN_188; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_190 = 6'h39 == io_index ? dirty_57 : _GEN_189; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_191 = 6'h3a == io_index ? dirty_58 : _GEN_190; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_192 = 6'h3b == io_index ? dirty_59 : _GEN_191; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_193 = 6'h3c == io_index ? dirty_60 : _GEN_192; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_194 = 6'h3d == io_index ? dirty_61 : _GEN_193; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_195 = 6'h3e == io_index ? dirty_62 : _GEN_194; // @[META.scala 31:24 META.scala 31:24]
  wire  _GEN_196 = 6'h3f == io_index ? dirty_63 : _GEN_195; // @[META.scala 31:24 META.scala 31:24]
  reg  io_valid_r_REG; // @[META.scala 32:24]
  wire  _GEN_198 = 6'h1 == io_index ? valid_1 : valid_0; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_199 = 6'h2 == io_index ? valid_2 : _GEN_198; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_200 = 6'h3 == io_index ? valid_3 : _GEN_199; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_201 = 6'h4 == io_index ? valid_4 : _GEN_200; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_202 = 6'h5 == io_index ? valid_5 : _GEN_201; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_203 = 6'h6 == io_index ? valid_6 : _GEN_202; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_204 = 6'h7 == io_index ? valid_7 : _GEN_203; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_205 = 6'h8 == io_index ? valid_8 : _GEN_204; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_206 = 6'h9 == io_index ? valid_9 : _GEN_205; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_207 = 6'ha == io_index ? valid_10 : _GEN_206; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_208 = 6'hb == io_index ? valid_11 : _GEN_207; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_209 = 6'hc == io_index ? valid_12 : _GEN_208; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_210 = 6'hd == io_index ? valid_13 : _GEN_209; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_211 = 6'he == io_index ? valid_14 : _GEN_210; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_212 = 6'hf == io_index ? valid_15 : _GEN_211; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_213 = 6'h10 == io_index ? valid_16 : _GEN_212; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_214 = 6'h11 == io_index ? valid_17 : _GEN_213; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_215 = 6'h12 == io_index ? valid_18 : _GEN_214; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_216 = 6'h13 == io_index ? valid_19 : _GEN_215; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_217 = 6'h14 == io_index ? valid_20 : _GEN_216; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_218 = 6'h15 == io_index ? valid_21 : _GEN_217; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_219 = 6'h16 == io_index ? valid_22 : _GEN_218; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_220 = 6'h17 == io_index ? valid_23 : _GEN_219; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_221 = 6'h18 == io_index ? valid_24 : _GEN_220; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_222 = 6'h19 == io_index ? valid_25 : _GEN_221; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_223 = 6'h1a == io_index ? valid_26 : _GEN_222; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_224 = 6'h1b == io_index ? valid_27 : _GEN_223; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_225 = 6'h1c == io_index ? valid_28 : _GEN_224; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_226 = 6'h1d == io_index ? valid_29 : _GEN_225; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_227 = 6'h1e == io_index ? valid_30 : _GEN_226; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_228 = 6'h1f == io_index ? valid_31 : _GEN_227; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_229 = 6'h20 == io_index ? valid_32 : _GEN_228; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_230 = 6'h21 == io_index ? valid_33 : _GEN_229; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_231 = 6'h22 == io_index ? valid_34 : _GEN_230; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_232 = 6'h23 == io_index ? valid_35 : _GEN_231; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_233 = 6'h24 == io_index ? valid_36 : _GEN_232; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_234 = 6'h25 == io_index ? valid_37 : _GEN_233; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_235 = 6'h26 == io_index ? valid_38 : _GEN_234; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_236 = 6'h27 == io_index ? valid_39 : _GEN_235; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_237 = 6'h28 == io_index ? valid_40 : _GEN_236; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_238 = 6'h29 == io_index ? valid_41 : _GEN_237; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_239 = 6'h2a == io_index ? valid_42 : _GEN_238; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_240 = 6'h2b == io_index ? valid_43 : _GEN_239; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_241 = 6'h2c == io_index ? valid_44 : _GEN_240; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_242 = 6'h2d == io_index ? valid_45 : _GEN_241; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_243 = 6'h2e == io_index ? valid_46 : _GEN_242; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_244 = 6'h2f == io_index ? valid_47 : _GEN_243; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_245 = 6'h30 == io_index ? valid_48 : _GEN_244; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_246 = 6'h31 == io_index ? valid_49 : _GEN_245; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_247 = 6'h32 == io_index ? valid_50 : _GEN_246; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_248 = 6'h33 == io_index ? valid_51 : _GEN_247; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_249 = 6'h34 == io_index ? valid_52 : _GEN_248; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_250 = 6'h35 == io_index ? valid_53 : _GEN_249; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_251 = 6'h36 == io_index ? valid_54 : _GEN_250; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_252 = 6'h37 == io_index ? valid_55 : _GEN_251; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_253 = 6'h38 == io_index ? valid_56 : _GEN_252; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_254 = 6'h39 == io_index ? valid_57 : _GEN_253; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_255 = 6'h3a == io_index ? valid_58 : _GEN_254; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_256 = 6'h3b == io_index ? valid_59 : _GEN_255; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_257 = 6'h3c == io_index ? valid_60 : _GEN_256; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_258 = 6'h3d == io_index ? valid_61 : _GEN_257; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_259 = 6'h3e == io_index ? valid_62 : _GEN_258; // @[META.scala 32:24 META.scala 32:24]
  wire  _GEN_260 = 6'h3f == io_index ? valid_63 : _GEN_259; // @[META.scala 32:24 META.scala 32:24]
  assign tag_io_tag_r_MPORT_addr = tag_io_tag_r_MPORT_addr_pipe_0;
  assign tag_io_tag_r_MPORT_data = tag[tag_io_tag_r_MPORT_addr]; // @[META.scala 20:24]
  assign tag_MPORT_data = io_tag_w;
  assign tag_MPORT_addr = io_index;
  assign tag_MPORT_mask = 1'h1;
  assign tag_MPORT_en = io_tag_wen;
  assign tag_MPORT_1_data = 22'h0;
  assign tag_MPORT_1_addr = 6'h0;
  assign tag_MPORT_1_mask = 1'h1;
  assign tag_MPORT_1_en = reset;
  assign tag_MPORT_2_data = 22'h0;
  assign tag_MPORT_2_addr = 6'h1;
  assign tag_MPORT_2_mask = 1'h1;
  assign tag_MPORT_2_en = reset;
  assign tag_MPORT_3_data = 22'h0;
  assign tag_MPORT_3_addr = 6'h2;
  assign tag_MPORT_3_mask = 1'h1;
  assign tag_MPORT_3_en = reset;
  assign tag_MPORT_4_data = 22'h0;
  assign tag_MPORT_4_addr = 6'h3;
  assign tag_MPORT_4_mask = 1'h1;
  assign tag_MPORT_4_en = reset;
  assign tag_MPORT_5_data = 22'h0;
  assign tag_MPORT_5_addr = 6'h4;
  assign tag_MPORT_5_mask = 1'h1;
  assign tag_MPORT_5_en = reset;
  assign tag_MPORT_6_data = 22'h0;
  assign tag_MPORT_6_addr = 6'h5;
  assign tag_MPORT_6_mask = 1'h1;
  assign tag_MPORT_6_en = reset;
  assign tag_MPORT_7_data = 22'h0;
  assign tag_MPORT_7_addr = 6'h6;
  assign tag_MPORT_7_mask = 1'h1;
  assign tag_MPORT_7_en = reset;
  assign tag_MPORT_8_data = 22'h0;
  assign tag_MPORT_8_addr = 6'h7;
  assign tag_MPORT_8_mask = 1'h1;
  assign tag_MPORT_8_en = reset;
  assign tag_MPORT_9_data = 22'h0;
  assign tag_MPORT_9_addr = 6'h8;
  assign tag_MPORT_9_mask = 1'h1;
  assign tag_MPORT_9_en = reset;
  assign tag_MPORT_10_data = 22'h0;
  assign tag_MPORT_10_addr = 6'h9;
  assign tag_MPORT_10_mask = 1'h1;
  assign tag_MPORT_10_en = reset;
  assign tag_MPORT_11_data = 22'h0;
  assign tag_MPORT_11_addr = 6'ha;
  assign tag_MPORT_11_mask = 1'h1;
  assign tag_MPORT_11_en = reset;
  assign tag_MPORT_12_data = 22'h0;
  assign tag_MPORT_12_addr = 6'hb;
  assign tag_MPORT_12_mask = 1'h1;
  assign tag_MPORT_12_en = reset;
  assign tag_MPORT_13_data = 22'h0;
  assign tag_MPORT_13_addr = 6'hc;
  assign tag_MPORT_13_mask = 1'h1;
  assign tag_MPORT_13_en = reset;
  assign tag_MPORT_14_data = 22'h0;
  assign tag_MPORT_14_addr = 6'hd;
  assign tag_MPORT_14_mask = 1'h1;
  assign tag_MPORT_14_en = reset;
  assign tag_MPORT_15_data = 22'h0;
  assign tag_MPORT_15_addr = 6'he;
  assign tag_MPORT_15_mask = 1'h1;
  assign tag_MPORT_15_en = reset;
  assign tag_MPORT_16_data = 22'h0;
  assign tag_MPORT_16_addr = 6'hf;
  assign tag_MPORT_16_mask = 1'h1;
  assign tag_MPORT_16_en = reset;
  assign tag_MPORT_17_data = 22'h0;
  assign tag_MPORT_17_addr = 6'h10;
  assign tag_MPORT_17_mask = 1'h1;
  assign tag_MPORT_17_en = reset;
  assign tag_MPORT_18_data = 22'h0;
  assign tag_MPORT_18_addr = 6'h11;
  assign tag_MPORT_18_mask = 1'h1;
  assign tag_MPORT_18_en = reset;
  assign tag_MPORT_19_data = 22'h0;
  assign tag_MPORT_19_addr = 6'h12;
  assign tag_MPORT_19_mask = 1'h1;
  assign tag_MPORT_19_en = reset;
  assign tag_MPORT_20_data = 22'h0;
  assign tag_MPORT_20_addr = 6'h13;
  assign tag_MPORT_20_mask = 1'h1;
  assign tag_MPORT_20_en = reset;
  assign tag_MPORT_21_data = 22'h0;
  assign tag_MPORT_21_addr = 6'h14;
  assign tag_MPORT_21_mask = 1'h1;
  assign tag_MPORT_21_en = reset;
  assign tag_MPORT_22_data = 22'h0;
  assign tag_MPORT_22_addr = 6'h15;
  assign tag_MPORT_22_mask = 1'h1;
  assign tag_MPORT_22_en = reset;
  assign tag_MPORT_23_data = 22'h0;
  assign tag_MPORT_23_addr = 6'h16;
  assign tag_MPORT_23_mask = 1'h1;
  assign tag_MPORT_23_en = reset;
  assign tag_MPORT_24_data = 22'h0;
  assign tag_MPORT_24_addr = 6'h17;
  assign tag_MPORT_24_mask = 1'h1;
  assign tag_MPORT_24_en = reset;
  assign tag_MPORT_25_data = 22'h0;
  assign tag_MPORT_25_addr = 6'h18;
  assign tag_MPORT_25_mask = 1'h1;
  assign tag_MPORT_25_en = reset;
  assign tag_MPORT_26_data = 22'h0;
  assign tag_MPORT_26_addr = 6'h19;
  assign tag_MPORT_26_mask = 1'h1;
  assign tag_MPORT_26_en = reset;
  assign tag_MPORT_27_data = 22'h0;
  assign tag_MPORT_27_addr = 6'h1a;
  assign tag_MPORT_27_mask = 1'h1;
  assign tag_MPORT_27_en = reset;
  assign tag_MPORT_28_data = 22'h0;
  assign tag_MPORT_28_addr = 6'h1b;
  assign tag_MPORT_28_mask = 1'h1;
  assign tag_MPORT_28_en = reset;
  assign tag_MPORT_29_data = 22'h0;
  assign tag_MPORT_29_addr = 6'h1c;
  assign tag_MPORT_29_mask = 1'h1;
  assign tag_MPORT_29_en = reset;
  assign tag_MPORT_30_data = 22'h0;
  assign tag_MPORT_30_addr = 6'h1d;
  assign tag_MPORT_30_mask = 1'h1;
  assign tag_MPORT_30_en = reset;
  assign tag_MPORT_31_data = 22'h0;
  assign tag_MPORT_31_addr = 6'h1e;
  assign tag_MPORT_31_mask = 1'h1;
  assign tag_MPORT_31_en = reset;
  assign tag_MPORT_32_data = 22'h0;
  assign tag_MPORT_32_addr = 6'h1f;
  assign tag_MPORT_32_mask = 1'h1;
  assign tag_MPORT_32_en = reset;
  assign tag_MPORT_33_data = 22'h0;
  assign tag_MPORT_33_addr = 6'h20;
  assign tag_MPORT_33_mask = 1'h1;
  assign tag_MPORT_33_en = reset;
  assign tag_MPORT_34_data = 22'h0;
  assign tag_MPORT_34_addr = 6'h21;
  assign tag_MPORT_34_mask = 1'h1;
  assign tag_MPORT_34_en = reset;
  assign tag_MPORT_35_data = 22'h0;
  assign tag_MPORT_35_addr = 6'h22;
  assign tag_MPORT_35_mask = 1'h1;
  assign tag_MPORT_35_en = reset;
  assign tag_MPORT_36_data = 22'h0;
  assign tag_MPORT_36_addr = 6'h23;
  assign tag_MPORT_36_mask = 1'h1;
  assign tag_MPORT_36_en = reset;
  assign tag_MPORT_37_data = 22'h0;
  assign tag_MPORT_37_addr = 6'h24;
  assign tag_MPORT_37_mask = 1'h1;
  assign tag_MPORT_37_en = reset;
  assign tag_MPORT_38_data = 22'h0;
  assign tag_MPORT_38_addr = 6'h25;
  assign tag_MPORT_38_mask = 1'h1;
  assign tag_MPORT_38_en = reset;
  assign tag_MPORT_39_data = 22'h0;
  assign tag_MPORT_39_addr = 6'h26;
  assign tag_MPORT_39_mask = 1'h1;
  assign tag_MPORT_39_en = reset;
  assign tag_MPORT_40_data = 22'h0;
  assign tag_MPORT_40_addr = 6'h27;
  assign tag_MPORT_40_mask = 1'h1;
  assign tag_MPORT_40_en = reset;
  assign tag_MPORT_41_data = 22'h0;
  assign tag_MPORT_41_addr = 6'h28;
  assign tag_MPORT_41_mask = 1'h1;
  assign tag_MPORT_41_en = reset;
  assign tag_MPORT_42_data = 22'h0;
  assign tag_MPORT_42_addr = 6'h29;
  assign tag_MPORT_42_mask = 1'h1;
  assign tag_MPORT_42_en = reset;
  assign tag_MPORT_43_data = 22'h0;
  assign tag_MPORT_43_addr = 6'h2a;
  assign tag_MPORT_43_mask = 1'h1;
  assign tag_MPORT_43_en = reset;
  assign tag_MPORT_44_data = 22'h0;
  assign tag_MPORT_44_addr = 6'h2b;
  assign tag_MPORT_44_mask = 1'h1;
  assign tag_MPORT_44_en = reset;
  assign tag_MPORT_45_data = 22'h0;
  assign tag_MPORT_45_addr = 6'h2c;
  assign tag_MPORT_45_mask = 1'h1;
  assign tag_MPORT_45_en = reset;
  assign tag_MPORT_46_data = 22'h0;
  assign tag_MPORT_46_addr = 6'h2d;
  assign tag_MPORT_46_mask = 1'h1;
  assign tag_MPORT_46_en = reset;
  assign tag_MPORT_47_data = 22'h0;
  assign tag_MPORT_47_addr = 6'h2e;
  assign tag_MPORT_47_mask = 1'h1;
  assign tag_MPORT_47_en = reset;
  assign tag_MPORT_48_data = 22'h0;
  assign tag_MPORT_48_addr = 6'h2f;
  assign tag_MPORT_48_mask = 1'h1;
  assign tag_MPORT_48_en = reset;
  assign tag_MPORT_49_data = 22'h0;
  assign tag_MPORT_49_addr = 6'h30;
  assign tag_MPORT_49_mask = 1'h1;
  assign tag_MPORT_49_en = reset;
  assign tag_MPORT_50_data = 22'h0;
  assign tag_MPORT_50_addr = 6'h31;
  assign tag_MPORT_50_mask = 1'h1;
  assign tag_MPORT_50_en = reset;
  assign tag_MPORT_51_data = 22'h0;
  assign tag_MPORT_51_addr = 6'h32;
  assign tag_MPORT_51_mask = 1'h1;
  assign tag_MPORT_51_en = reset;
  assign tag_MPORT_52_data = 22'h0;
  assign tag_MPORT_52_addr = 6'h33;
  assign tag_MPORT_52_mask = 1'h1;
  assign tag_MPORT_52_en = reset;
  assign tag_MPORT_53_data = 22'h0;
  assign tag_MPORT_53_addr = 6'h34;
  assign tag_MPORT_53_mask = 1'h1;
  assign tag_MPORT_53_en = reset;
  assign tag_MPORT_54_data = 22'h0;
  assign tag_MPORT_54_addr = 6'h35;
  assign tag_MPORT_54_mask = 1'h1;
  assign tag_MPORT_54_en = reset;
  assign tag_MPORT_55_data = 22'h0;
  assign tag_MPORT_55_addr = 6'h36;
  assign tag_MPORT_55_mask = 1'h1;
  assign tag_MPORT_55_en = reset;
  assign tag_MPORT_56_data = 22'h0;
  assign tag_MPORT_56_addr = 6'h37;
  assign tag_MPORT_56_mask = 1'h1;
  assign tag_MPORT_56_en = reset;
  assign tag_MPORT_57_data = 22'h0;
  assign tag_MPORT_57_addr = 6'h38;
  assign tag_MPORT_57_mask = 1'h1;
  assign tag_MPORT_57_en = reset;
  assign tag_MPORT_58_data = 22'h0;
  assign tag_MPORT_58_addr = 6'h39;
  assign tag_MPORT_58_mask = 1'h1;
  assign tag_MPORT_58_en = reset;
  assign tag_MPORT_59_data = 22'h0;
  assign tag_MPORT_59_addr = 6'h3a;
  assign tag_MPORT_59_mask = 1'h1;
  assign tag_MPORT_59_en = reset;
  assign tag_MPORT_60_data = 22'h0;
  assign tag_MPORT_60_addr = 6'h3b;
  assign tag_MPORT_60_mask = 1'h1;
  assign tag_MPORT_60_en = reset;
  assign tag_MPORT_61_data = 22'h0;
  assign tag_MPORT_61_addr = 6'h3c;
  assign tag_MPORT_61_mask = 1'h1;
  assign tag_MPORT_61_en = reset;
  assign tag_MPORT_62_data = 22'h0;
  assign tag_MPORT_62_addr = 6'h3d;
  assign tag_MPORT_62_mask = 1'h1;
  assign tag_MPORT_62_en = reset;
  assign tag_MPORT_63_data = 22'h0;
  assign tag_MPORT_63_addr = 6'h3e;
  assign tag_MPORT_63_mask = 1'h1;
  assign tag_MPORT_63_en = reset;
  assign tag_MPORT_64_data = 22'h0;
  assign tag_MPORT_64_addr = 6'h3f;
  assign tag_MPORT_64_mask = 1'h1;
  assign tag_MPORT_64_en = reset;
  assign io_tag_r = tag_io_tag_r_MPORT_data; // @[META.scala 29:12]
  assign io_dirty_r = io_dirty_r_REG; // @[META.scala 31:14]
  assign io_valid_r = io_valid_r_REG; // @[META.scala 32:14]
  assign io_fence_dirty = _GEN_196 & _GEN_260; // @[META.scala 33:34]
  always @(posedge clock) begin
    if(tag_MPORT_en & tag_MPORT_mask) begin
      tag[tag_MPORT_addr] <= tag_MPORT_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_1_en & tag_MPORT_1_mask) begin
      tag[tag_MPORT_1_addr] <= tag_MPORT_1_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_2_en & tag_MPORT_2_mask) begin
      tag[tag_MPORT_2_addr] <= tag_MPORT_2_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_3_en & tag_MPORT_3_mask) begin
      tag[tag_MPORT_3_addr] <= tag_MPORT_3_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_4_en & tag_MPORT_4_mask) begin
      tag[tag_MPORT_4_addr] <= tag_MPORT_4_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_5_en & tag_MPORT_5_mask) begin
      tag[tag_MPORT_5_addr] <= tag_MPORT_5_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_6_en & tag_MPORT_6_mask) begin
      tag[tag_MPORT_6_addr] <= tag_MPORT_6_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_7_en & tag_MPORT_7_mask) begin
      tag[tag_MPORT_7_addr] <= tag_MPORT_7_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_8_en & tag_MPORT_8_mask) begin
      tag[tag_MPORT_8_addr] <= tag_MPORT_8_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_9_en & tag_MPORT_9_mask) begin
      tag[tag_MPORT_9_addr] <= tag_MPORT_9_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_10_en & tag_MPORT_10_mask) begin
      tag[tag_MPORT_10_addr] <= tag_MPORT_10_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_11_en & tag_MPORT_11_mask) begin
      tag[tag_MPORT_11_addr] <= tag_MPORT_11_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_12_en & tag_MPORT_12_mask) begin
      tag[tag_MPORT_12_addr] <= tag_MPORT_12_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_13_en & tag_MPORT_13_mask) begin
      tag[tag_MPORT_13_addr] <= tag_MPORT_13_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_14_en & tag_MPORT_14_mask) begin
      tag[tag_MPORT_14_addr] <= tag_MPORT_14_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_15_en & tag_MPORT_15_mask) begin
      tag[tag_MPORT_15_addr] <= tag_MPORT_15_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_16_en & tag_MPORT_16_mask) begin
      tag[tag_MPORT_16_addr] <= tag_MPORT_16_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_17_en & tag_MPORT_17_mask) begin
      tag[tag_MPORT_17_addr] <= tag_MPORT_17_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_18_en & tag_MPORT_18_mask) begin
      tag[tag_MPORT_18_addr] <= tag_MPORT_18_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_19_en & tag_MPORT_19_mask) begin
      tag[tag_MPORT_19_addr] <= tag_MPORT_19_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_20_en & tag_MPORT_20_mask) begin
      tag[tag_MPORT_20_addr] <= tag_MPORT_20_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_21_en & tag_MPORT_21_mask) begin
      tag[tag_MPORT_21_addr] <= tag_MPORT_21_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_22_en & tag_MPORT_22_mask) begin
      tag[tag_MPORT_22_addr] <= tag_MPORT_22_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_23_en & tag_MPORT_23_mask) begin
      tag[tag_MPORT_23_addr] <= tag_MPORT_23_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_24_en & tag_MPORT_24_mask) begin
      tag[tag_MPORT_24_addr] <= tag_MPORT_24_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_25_en & tag_MPORT_25_mask) begin
      tag[tag_MPORT_25_addr] <= tag_MPORT_25_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_26_en & tag_MPORT_26_mask) begin
      tag[tag_MPORT_26_addr] <= tag_MPORT_26_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_27_en & tag_MPORT_27_mask) begin
      tag[tag_MPORT_27_addr] <= tag_MPORT_27_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_28_en & tag_MPORT_28_mask) begin
      tag[tag_MPORT_28_addr] <= tag_MPORT_28_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_29_en & tag_MPORT_29_mask) begin
      tag[tag_MPORT_29_addr] <= tag_MPORT_29_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_30_en & tag_MPORT_30_mask) begin
      tag[tag_MPORT_30_addr] <= tag_MPORT_30_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_31_en & tag_MPORT_31_mask) begin
      tag[tag_MPORT_31_addr] <= tag_MPORT_31_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_32_en & tag_MPORT_32_mask) begin
      tag[tag_MPORT_32_addr] <= tag_MPORT_32_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_33_en & tag_MPORT_33_mask) begin
      tag[tag_MPORT_33_addr] <= tag_MPORT_33_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_34_en & tag_MPORT_34_mask) begin
      tag[tag_MPORT_34_addr] <= tag_MPORT_34_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_35_en & tag_MPORT_35_mask) begin
      tag[tag_MPORT_35_addr] <= tag_MPORT_35_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_36_en & tag_MPORT_36_mask) begin
      tag[tag_MPORT_36_addr] <= tag_MPORT_36_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_37_en & tag_MPORT_37_mask) begin
      tag[tag_MPORT_37_addr] <= tag_MPORT_37_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_38_en & tag_MPORT_38_mask) begin
      tag[tag_MPORT_38_addr] <= tag_MPORT_38_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_39_en & tag_MPORT_39_mask) begin
      tag[tag_MPORT_39_addr] <= tag_MPORT_39_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_40_en & tag_MPORT_40_mask) begin
      tag[tag_MPORT_40_addr] <= tag_MPORT_40_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_41_en & tag_MPORT_41_mask) begin
      tag[tag_MPORT_41_addr] <= tag_MPORT_41_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_42_en & tag_MPORT_42_mask) begin
      tag[tag_MPORT_42_addr] <= tag_MPORT_42_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_43_en & tag_MPORT_43_mask) begin
      tag[tag_MPORT_43_addr] <= tag_MPORT_43_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_44_en & tag_MPORT_44_mask) begin
      tag[tag_MPORT_44_addr] <= tag_MPORT_44_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_45_en & tag_MPORT_45_mask) begin
      tag[tag_MPORT_45_addr] <= tag_MPORT_45_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_46_en & tag_MPORT_46_mask) begin
      tag[tag_MPORT_46_addr] <= tag_MPORT_46_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_47_en & tag_MPORT_47_mask) begin
      tag[tag_MPORT_47_addr] <= tag_MPORT_47_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_48_en & tag_MPORT_48_mask) begin
      tag[tag_MPORT_48_addr] <= tag_MPORT_48_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_49_en & tag_MPORT_49_mask) begin
      tag[tag_MPORT_49_addr] <= tag_MPORT_49_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_50_en & tag_MPORT_50_mask) begin
      tag[tag_MPORT_50_addr] <= tag_MPORT_50_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_51_en & tag_MPORT_51_mask) begin
      tag[tag_MPORT_51_addr] <= tag_MPORT_51_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_52_en & tag_MPORT_52_mask) begin
      tag[tag_MPORT_52_addr] <= tag_MPORT_52_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_53_en & tag_MPORT_53_mask) begin
      tag[tag_MPORT_53_addr] <= tag_MPORT_53_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_54_en & tag_MPORT_54_mask) begin
      tag[tag_MPORT_54_addr] <= tag_MPORT_54_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_55_en & tag_MPORT_55_mask) begin
      tag[tag_MPORT_55_addr] <= tag_MPORT_55_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_56_en & tag_MPORT_56_mask) begin
      tag[tag_MPORT_56_addr] <= tag_MPORT_56_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_57_en & tag_MPORT_57_mask) begin
      tag[tag_MPORT_57_addr] <= tag_MPORT_57_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_58_en & tag_MPORT_58_mask) begin
      tag[tag_MPORT_58_addr] <= tag_MPORT_58_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_59_en & tag_MPORT_59_mask) begin
      tag[tag_MPORT_59_addr] <= tag_MPORT_59_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_60_en & tag_MPORT_60_mask) begin
      tag[tag_MPORT_60_addr] <= tag_MPORT_60_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_61_en & tag_MPORT_61_mask) begin
      tag[tag_MPORT_61_addr] <= tag_MPORT_61_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_62_en & tag_MPORT_62_mask) begin
      tag[tag_MPORT_62_addr] <= tag_MPORT_62_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_63_en & tag_MPORT_63_mask) begin
      tag[tag_MPORT_63_addr] <= tag_MPORT_63_data; // @[META.scala 20:24]
    end
    if(tag_MPORT_64_en & tag_MPORT_64_mask) begin
      tag[tag_MPORT_64_addr] <= tag_MPORT_64_data; // @[META.scala 20:24]
    end
    tag_io_tag_r_MPORT_addr_pipe_0 <= io_index;
    if (reset) begin // @[META.scala 22:22]
      valid_0 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_0 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_0 <= _GEN_0;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_1 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_1 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_1 <= _GEN_1;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_2 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_2 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_2 <= _GEN_2;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_3 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_3 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_3 <= _GEN_3;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_4 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_4 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_4 <= _GEN_4;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_5 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_5 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_5 <= _GEN_5;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_6 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_6 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_6 <= _GEN_6;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_7 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_7 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_7 <= _GEN_7;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_8 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_8 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_8 <= _GEN_8;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_9 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_9 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_9 <= _GEN_9;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_10 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_10 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_10 <= _GEN_10;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_11 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_11 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_11 <= _GEN_11;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_12 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_12 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_12 <= _GEN_12;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_13 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_13 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_13 <= _GEN_13;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_14 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_14 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_14 <= _GEN_14;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_15 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_15 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_15 <= _GEN_15;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_16 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_16 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_16 <= _GEN_16;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_17 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_17 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_17 <= _GEN_17;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_18 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_18 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_18 <= _GEN_18;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_19 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_19 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_19 <= _GEN_19;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_20 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_20 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_20 <= _GEN_20;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_21 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_21 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_21 <= _GEN_21;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_22 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_22 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_22 <= _GEN_22;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_23 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_23 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_23 <= _GEN_23;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_24 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_24 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_24 <= _GEN_24;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_25 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_25 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_25 <= _GEN_25;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_26 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_26 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_26 <= _GEN_26;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_27 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_27 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_27 <= _GEN_27;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_28 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_28 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_28 <= _GEN_28;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_29 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_29 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_29 <= _GEN_29;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_30 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_30 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_30 <= _GEN_30;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_31 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_31 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_31 <= _GEN_31;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_32 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_32 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_32 <= _GEN_32;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_33 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_33 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_33 <= _GEN_33;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_34 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_34 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_34 <= _GEN_34;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_35 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_35 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_35 <= _GEN_35;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_36 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_36 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_36 <= _GEN_36;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_37 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_37 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_37 <= _GEN_37;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_38 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_38 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_38 <= _GEN_38;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_39 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_39 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_39 <= _GEN_39;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_40 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_40 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_40 <= _GEN_40;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_41 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_41 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_41 <= _GEN_41;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_42 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_42 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_42 <= _GEN_42;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_43 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_43 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_43 <= _GEN_43;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_44 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_44 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_44 <= _GEN_44;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_45 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_45 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_45 <= _GEN_45;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_46 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_46 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_46 <= _GEN_46;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_47 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_47 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_47 <= _GEN_47;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_48 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_48 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_48 <= _GEN_48;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_49 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_49 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_49 <= _GEN_49;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_50 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_50 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_50 <= _GEN_50;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_51 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_51 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_51 <= _GEN_51;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_52 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_52 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_52 <= _GEN_52;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_53 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_53 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_53 <= _GEN_53;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_54 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_54 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_54 <= _GEN_54;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_55 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_55 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_55 <= _GEN_55;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_56 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_56 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_56 <= _GEN_56;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_57 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_57 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_57 <= _GEN_57;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_58 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_58 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_58 <= _GEN_58;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_59 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_59 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_59 <= _GEN_59;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_60 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_60 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_60 <= _GEN_60;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_61 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_61 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_61 <= _GEN_61;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_62 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_62 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_62 <= _GEN_62;
    end
    if (reset) begin // @[META.scala 22:22]
      valid_63 <= 1'h0; // @[META.scala 22:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      valid_63 <= 1'h0; // @[META.scala 48:16]
    end else if (io_tag_wen) begin // @[META.scala 25:21]
      valid_63 <= _GEN_63;
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_0 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_0 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h0 == io_index) begin // @[META.scala 36:18]
        dirty_0 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_1 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_1 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1 == io_index) begin // @[META.scala 36:18]
        dirty_1 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_2 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_2 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2 == io_index) begin // @[META.scala 36:18]
        dirty_2 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_3 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_3 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3 == io_index) begin // @[META.scala 36:18]
        dirty_3 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_4 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_4 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h4 == io_index) begin // @[META.scala 36:18]
        dirty_4 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_5 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_5 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h5 == io_index) begin // @[META.scala 36:18]
        dirty_5 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_6 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_6 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h6 == io_index) begin // @[META.scala 36:18]
        dirty_6 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_7 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_7 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h7 == io_index) begin // @[META.scala 36:18]
        dirty_7 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_8 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_8 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h8 == io_index) begin // @[META.scala 36:18]
        dirty_8 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_9 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_9 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h9 == io_index) begin // @[META.scala 36:18]
        dirty_9 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_10 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_10 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'ha == io_index) begin // @[META.scala 36:18]
        dirty_10 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_11 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_11 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'hb == io_index) begin // @[META.scala 36:18]
        dirty_11 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_12 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_12 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'hc == io_index) begin // @[META.scala 36:18]
        dirty_12 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_13 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_13 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'hd == io_index) begin // @[META.scala 36:18]
        dirty_13 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_14 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_14 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'he == io_index) begin // @[META.scala 36:18]
        dirty_14 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_15 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_15 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'hf == io_index) begin // @[META.scala 36:18]
        dirty_15 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_16 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_16 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h10 == io_index) begin // @[META.scala 36:18]
        dirty_16 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_17 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_17 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h11 == io_index) begin // @[META.scala 36:18]
        dirty_17 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_18 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_18 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h12 == io_index) begin // @[META.scala 36:18]
        dirty_18 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_19 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_19 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h13 == io_index) begin // @[META.scala 36:18]
        dirty_19 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_20 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_20 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h14 == io_index) begin // @[META.scala 36:18]
        dirty_20 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_21 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_21 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h15 == io_index) begin // @[META.scala 36:18]
        dirty_21 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_22 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_22 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h16 == io_index) begin // @[META.scala 36:18]
        dirty_22 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_23 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_23 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h17 == io_index) begin // @[META.scala 36:18]
        dirty_23 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_24 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_24 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h18 == io_index) begin // @[META.scala 36:18]
        dirty_24 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_25 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_25 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h19 == io_index) begin // @[META.scala 36:18]
        dirty_25 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_26 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_26 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1a == io_index) begin // @[META.scala 36:18]
        dirty_26 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_27 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_27 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1b == io_index) begin // @[META.scala 36:18]
        dirty_27 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_28 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_28 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1c == io_index) begin // @[META.scala 36:18]
        dirty_28 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_29 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_29 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1d == io_index) begin // @[META.scala 36:18]
        dirty_29 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_30 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_30 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1e == io_index) begin // @[META.scala 36:18]
        dirty_30 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_31 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_31 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h1f == io_index) begin // @[META.scala 36:18]
        dirty_31 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_32 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_32 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h20 == io_index) begin // @[META.scala 36:18]
        dirty_32 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_33 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_33 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h21 == io_index) begin // @[META.scala 36:18]
        dirty_33 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_34 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_34 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h22 == io_index) begin // @[META.scala 36:18]
        dirty_34 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_35 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_35 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h23 == io_index) begin // @[META.scala 36:18]
        dirty_35 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_36 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_36 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h24 == io_index) begin // @[META.scala 36:18]
        dirty_36 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_37 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_37 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h25 == io_index) begin // @[META.scala 36:18]
        dirty_37 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_38 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_38 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h26 == io_index) begin // @[META.scala 36:18]
        dirty_38 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_39 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_39 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h27 == io_index) begin // @[META.scala 36:18]
        dirty_39 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_40 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_40 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h28 == io_index) begin // @[META.scala 36:18]
        dirty_40 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_41 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_41 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h29 == io_index) begin // @[META.scala 36:18]
        dirty_41 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_42 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_42 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2a == io_index) begin // @[META.scala 36:18]
        dirty_42 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_43 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_43 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2b == io_index) begin // @[META.scala 36:18]
        dirty_43 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_44 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_44 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2c == io_index) begin // @[META.scala 36:18]
        dirty_44 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_45 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_45 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2d == io_index) begin // @[META.scala 36:18]
        dirty_45 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_46 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_46 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2e == io_index) begin // @[META.scala 36:18]
        dirty_46 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_47 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_47 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h2f == io_index) begin // @[META.scala 36:18]
        dirty_47 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_48 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_48 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h30 == io_index) begin // @[META.scala 36:18]
        dirty_48 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_49 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_49 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h31 == io_index) begin // @[META.scala 36:18]
        dirty_49 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_50 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_50 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h32 == io_index) begin // @[META.scala 36:18]
        dirty_50 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_51 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_51 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h33 == io_index) begin // @[META.scala 36:18]
        dirty_51 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_52 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_52 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h34 == io_index) begin // @[META.scala 36:18]
        dirty_52 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_53 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_53 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h35 == io_index) begin // @[META.scala 36:18]
        dirty_53 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_54 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_54 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h36 == io_index) begin // @[META.scala 36:18]
        dirty_54 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_55 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_55 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h37 == io_index) begin // @[META.scala 36:18]
        dirty_55 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_56 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_56 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h38 == io_index) begin // @[META.scala 36:18]
        dirty_56 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_57 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_57 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h39 == io_index) begin // @[META.scala 36:18]
        dirty_57 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_58 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_58 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3a == io_index) begin // @[META.scala 36:18]
        dirty_58 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_59 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_59 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3b == io_index) begin // @[META.scala 36:18]
        dirty_59 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_60 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_60 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3c == io_index) begin // @[META.scala 36:18]
        dirty_60 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_61 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_61 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3d == io_index) begin // @[META.scala 36:18]
        dirty_61 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_62 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_62 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3e == io_index) begin // @[META.scala 36:18]
        dirty_62 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 23:22]
      dirty_63 <= 1'h0; // @[META.scala 23:22]
    end else if (io_fence) begin // @[META.scala 45:19]
      dirty_63 <= 1'h0; // @[META.scala 47:16]
    end else if (io_dirty_wen) begin // @[META.scala 35:23]
      if (6'h3f == io_index) begin // @[META.scala 36:18]
        dirty_63 <= io_dirty_w; // @[META.scala 36:18]
      end
    end
    if (reset) begin // @[META.scala 31:24]
      io_dirty_r_REG <= 1'h0; // @[META.scala 31:24]
    end else if (6'h3f == io_index) begin // @[META.scala 31:24]
      io_dirty_r_REG <= dirty_63; // @[META.scala 31:24]
    end else if (6'h3e == io_index) begin // @[META.scala 31:24]
      io_dirty_r_REG <= dirty_62; // @[META.scala 31:24]
    end else if (6'h3d == io_index) begin // @[META.scala 31:24]
      io_dirty_r_REG <= dirty_61; // @[META.scala 31:24]
    end else begin
      io_dirty_r_REG <= _GEN_193;
    end
    if (reset) begin // @[META.scala 32:24]
      io_valid_r_REG <= 1'h0; // @[META.scala 32:24]
    end else if (6'h3f == io_index) begin // @[META.scala 32:24]
      io_valid_r_REG <= valid_63; // @[META.scala 32:24]
    end else if (6'h3e == io_index) begin // @[META.scala 32:24]
      io_valid_r_REG <= valid_62; // @[META.scala 32:24]
    end else if (6'h3d == io_index) begin // @[META.scala 32:24]
      io_valid_r_REG <= valid_61; // @[META.scala 32:24]
    end else begin
      io_valid_r_REG <= _GEN_257;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag[initvar] = _RAND_0[21:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tag_io_tag_r_MPORT_addr_pipe_0 = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  valid_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_3 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_4 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_5 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_6 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_7 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_8 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_9 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_10 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_11 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_12 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_13 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_14 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_15 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_16 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_17 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_18 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_19 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_20 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_21 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_22 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_23 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_24 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_25 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_26 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_27 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_28 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_29 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_30 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_31 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_32 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_33 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_34 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_35 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_36 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_37 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_38 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_39 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_40 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_41 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_42 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_43 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_44 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_45 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_46 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_47 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_48 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_49 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_50 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_51 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_52 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_53 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_54 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_55 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_56 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_57 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_58 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_59 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_60 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_61 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_62 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_63 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  dirty_0 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  dirty_1 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  dirty_2 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  dirty_3 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  dirty_4 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  dirty_5 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  dirty_6 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  dirty_7 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  dirty_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  dirty_9 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  dirty_10 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  dirty_11 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  dirty_12 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  dirty_13 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  dirty_14 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  dirty_15 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  dirty_16 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  dirty_17 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  dirty_18 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  dirty_19 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  dirty_20 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  dirty_21 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  dirty_22 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  dirty_23 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  dirty_24 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  dirty_25 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  dirty_26 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  dirty_27 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  dirty_28 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  dirty_29 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  dirty_30 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  dirty_31 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  dirty_32 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  dirty_33 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  dirty_34 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  dirty_35 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  dirty_36 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  dirty_37 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  dirty_38 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  dirty_39 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  dirty_40 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  dirty_41 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  dirty_42 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  dirty_43 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  dirty_44 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  dirty_45 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  dirty_46 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  dirty_47 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  dirty_48 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  dirty_49 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  dirty_50 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  dirty_51 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  dirty_52 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  dirty_53 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  dirty_54 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  dirty_55 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  dirty_56 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  dirty_57 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  dirty_58 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  dirty_59 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  dirty_60 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  dirty_61 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  dirty_62 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  dirty_63 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  io_dirty_r_REG = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  io_valid_r_REG = _RAND_131[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Cache_Soc(
  input          clock,
  input          reset,
  input          io_in_valid,
  input          io_in_op,
  input  [31:0]  io_in_addr,
  input  [7:0]   io_in_wstrb,
  input  [63:0]  io_in_wdata,
  input          io_in_fence,
  output         io_in_fence_finish,
  output         io_in_data_ok,
  output [63:0]  io_in_rdata,
  output [127:0] io_in_inst,
  output         io_out_rd_req,
  output [2:0]   io_out_rd_size,
  output [31:0]  io_out_rd_addr,
  input          io_out_rd_rdy,
  input          io_out_ret_valid,
  input  [127:0] io_out_ret_data,
  output         io_out_wr_req,
  output [2:0]   io_out_wr_size,
  output [31:0]  io_out_wr_addr,
  output [7:0]   io_out_wr_wstrb,
  output [127:0] io_out_wr_data,
  input          io_out_wr_rdy,
  input          io_out_wr_ok,
  output         io_sram_0_en,
  output         io_sram_0_wen,
  output [5:0]   io_sram_0_addr,
  output [127:0] io_sram_0_wdata,
  input  [127:0] io_sram_0_rdata,
  output         io_sram_1_en,
  output         io_sram_1_wen,
  output [5:0]   io_sram_1_addr,
  output [127:0] io_sram_1_wdata,
  input  [127:0] io_sram_1_rdata,
  output         io_sram_2_en,
  output         io_sram_2_wen,
  output [5:0]   io_sram_2_addr,
  output [127:0] io_sram_2_wdata,
  input  [127:0] io_sram_2_rdata,
  output         io_sram_3_en,
  output         io_sram_3_wen,
  output [5:0]   io_sram_3_addr,
  output [127:0] io_sram_3_wdata,
  input  [127:0] io_sram_3_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
`endif // RANDOMIZE_REG_INIT
  wire  meta_0_clock; // @[Cache_Soc.scala 24:22]
  wire  meta_0_reset; // @[Cache_Soc.scala 24:22]
  wire [5:0] meta_0_io_index; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_0_io_tag_r; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_0_io_tag_w; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_tag_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_dirty_r; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_dirty_w; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_dirty_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_valid_r; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_fence; // @[Cache_Soc.scala 24:22]
  wire  meta_0_io_fence_dirty; // @[Cache_Soc.scala 24:22]
  wire  meta_1_clock; // @[Cache_Soc.scala 24:22]
  wire  meta_1_reset; // @[Cache_Soc.scala 24:22]
  wire [5:0] meta_1_io_index; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_1_io_tag_r; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_1_io_tag_w; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_tag_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_dirty_r; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_dirty_w; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_dirty_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_valid_r; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_fence; // @[Cache_Soc.scala 24:22]
  wire  meta_1_io_fence_dirty; // @[Cache_Soc.scala 24:22]
  wire  meta_2_clock; // @[Cache_Soc.scala 24:22]
  wire  meta_2_reset; // @[Cache_Soc.scala 24:22]
  wire [5:0] meta_2_io_index; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_2_io_tag_r; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_2_io_tag_w; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_tag_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_dirty_r; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_dirty_w; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_dirty_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_valid_r; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_fence; // @[Cache_Soc.scala 24:22]
  wire  meta_2_io_fence_dirty; // @[Cache_Soc.scala 24:22]
  wire  meta_3_clock; // @[Cache_Soc.scala 24:22]
  wire  meta_3_reset; // @[Cache_Soc.scala 24:22]
  wire [5:0] meta_3_io_index; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_3_io_tag_r; // @[Cache_Soc.scala 24:22]
  wire [21:0] meta_3_io_tag_w; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_tag_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_dirty_r; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_dirty_w; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_dirty_wen; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_valid_r; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_fence; // @[Cache_Soc.scala 24:22]
  wire  meta_3_io_fence_dirty; // @[Cache_Soc.scala 24:22]
  reg [2:0] state; // @[Cache_Soc.scala 41:22]
  reg  wb_state; // @[Cache_Soc.scala 42:25]
  reg [2:0] fence_state; // @[Cache_Soc.scala 43:28]
  wire  in_uncache = ~io_in_addr[31]; // @[Cache_Soc.scala 49:20]
  wire [5:0] in_index = io_in_addr[9:4]; // @[Cache_Soc.scala 50:25]
  wire [21:0] in_tag = io_in_addr[31:10]; // @[Cache_Soc.scala 51:23]
  wire [3:0] in_offset = io_in_addr[3:0]; // @[Cache_Soc.scala 52:26]
  reg  rb_op; // @[Cache_Soc.scala 55:22]
  reg  rb_uncache; // @[Cache_Soc.scala 56:27]
  reg [5:0] rb_index; // @[Cache_Soc.scala 57:25]
  reg [21:0] rb_tag; // @[Cache_Soc.scala 58:23]
  reg [3:0] rb_offset; // @[Cache_Soc.scala 59:26]
  reg [7:0] rb_wstrb; // @[Cache_Soc.scala 60:25]
  reg [63:0] rb_wdata; // @[Cache_Soc.scala 61:25]
  reg [1:0] wb_hitway; // @[Cache_Soc.scala 64:26]
  reg [5:0] wb_index; // @[Cache_Soc.scala 65:25]
  reg [3:0] wb_offset; // @[Cache_Soc.scala 67:26]
  reg [7:0] wb_wstrb; // @[Cache_Soc.scala 68:25]
  reg [63:0] wb_wdata; // @[Cache_Soc.scala 69:25]
  reg  replace_valid; // @[Cache_Soc.scala 72:30]
  reg  replace_dirty; // @[Cache_Soc.scala 73:30]
  reg [21:0] replace_tag; // @[Cache_Soc.scala 74:28]
  reg [127:0] replace_data; // @[Cache_Soc.scala 75:29]
  wire [21:0] tag_0 = meta_0_io_tag_r;
  wire  valid_0 = meta_0_io_valid_r;
  wire  hit_0 = tag_0 == rb_tag & valid_0; // @[Cache_Soc.scala 85:25]
  wire [21:0] tag_1 = meta_1_io_tag_r;
  wire  valid_1 = meta_1_io_valid_r;
  wire  hit_1 = tag_1 == rb_tag & valid_1; // @[Cache_Soc.scala 85:25]
  wire [21:0] tag_2 = meta_2_io_tag_r;
  wire  valid_2 = meta_2_io_valid_r;
  wire  hit_2 = tag_2 == rb_tag & valid_2; // @[Cache_Soc.scala 85:25]
  wire [21:0] tag_3 = meta_3_io_tag_r;
  wire  valid_3 = meta_3_io_valid_r;
  wire  hit_3 = tag_3 == rb_tag & valid_3; // @[Cache_Soc.scala 85:25]
  wire [3:0] _cache_hit_T = {hit_0,hit_1,hit_2,hit_3}; // @[Cat.scala 30:58]
  wire  _cache_hit_T_2 = ~rb_uncache; // @[Cache_Soc.scala 87:32]
  wire  cache_hit = |_cache_hit_T & ~rb_uncache; // @[Cache_Soc.scala 87:29]
  reg  plru0_0; // @[Cache_Soc.scala 89:22]
  reg  plru0_1; // @[Cache_Soc.scala 89:22]
  reg  plru0_2; // @[Cache_Soc.scala 89:22]
  reg  plru0_3; // @[Cache_Soc.scala 89:22]
  reg  plru0_4; // @[Cache_Soc.scala 89:22]
  reg  plru0_5; // @[Cache_Soc.scala 89:22]
  reg  plru0_6; // @[Cache_Soc.scala 89:22]
  reg  plru0_7; // @[Cache_Soc.scala 89:22]
  reg  plru0_8; // @[Cache_Soc.scala 89:22]
  reg  plru0_9; // @[Cache_Soc.scala 89:22]
  reg  plru0_10; // @[Cache_Soc.scala 89:22]
  reg  plru0_11; // @[Cache_Soc.scala 89:22]
  reg  plru0_12; // @[Cache_Soc.scala 89:22]
  reg  plru0_13; // @[Cache_Soc.scala 89:22]
  reg  plru0_14; // @[Cache_Soc.scala 89:22]
  reg  plru0_15; // @[Cache_Soc.scala 89:22]
  reg  plru0_16; // @[Cache_Soc.scala 89:22]
  reg  plru0_17; // @[Cache_Soc.scala 89:22]
  reg  plru0_18; // @[Cache_Soc.scala 89:22]
  reg  plru0_19; // @[Cache_Soc.scala 89:22]
  reg  plru0_20; // @[Cache_Soc.scala 89:22]
  reg  plru0_21; // @[Cache_Soc.scala 89:22]
  reg  plru0_22; // @[Cache_Soc.scala 89:22]
  reg  plru0_23; // @[Cache_Soc.scala 89:22]
  reg  plru0_24; // @[Cache_Soc.scala 89:22]
  reg  plru0_25; // @[Cache_Soc.scala 89:22]
  reg  plru0_26; // @[Cache_Soc.scala 89:22]
  reg  plru0_27; // @[Cache_Soc.scala 89:22]
  reg  plru0_28; // @[Cache_Soc.scala 89:22]
  reg  plru0_29; // @[Cache_Soc.scala 89:22]
  reg  plru0_30; // @[Cache_Soc.scala 89:22]
  reg  plru0_31; // @[Cache_Soc.scala 89:22]
  reg  plru0_32; // @[Cache_Soc.scala 89:22]
  reg  plru0_33; // @[Cache_Soc.scala 89:22]
  reg  plru0_34; // @[Cache_Soc.scala 89:22]
  reg  plru0_35; // @[Cache_Soc.scala 89:22]
  reg  plru0_36; // @[Cache_Soc.scala 89:22]
  reg  plru0_37; // @[Cache_Soc.scala 89:22]
  reg  plru0_38; // @[Cache_Soc.scala 89:22]
  reg  plru0_39; // @[Cache_Soc.scala 89:22]
  reg  plru0_40; // @[Cache_Soc.scala 89:22]
  reg  plru0_41; // @[Cache_Soc.scala 89:22]
  reg  plru0_42; // @[Cache_Soc.scala 89:22]
  reg  plru0_43; // @[Cache_Soc.scala 89:22]
  reg  plru0_44; // @[Cache_Soc.scala 89:22]
  reg  plru0_45; // @[Cache_Soc.scala 89:22]
  reg  plru0_46; // @[Cache_Soc.scala 89:22]
  reg  plru0_47; // @[Cache_Soc.scala 89:22]
  reg  plru0_48; // @[Cache_Soc.scala 89:22]
  reg  plru0_49; // @[Cache_Soc.scala 89:22]
  reg  plru0_50; // @[Cache_Soc.scala 89:22]
  reg  plru0_51; // @[Cache_Soc.scala 89:22]
  reg  plru0_52; // @[Cache_Soc.scala 89:22]
  reg  plru0_53; // @[Cache_Soc.scala 89:22]
  reg  plru0_54; // @[Cache_Soc.scala 89:22]
  reg  plru0_55; // @[Cache_Soc.scala 89:22]
  reg  plru0_56; // @[Cache_Soc.scala 89:22]
  reg  plru0_57; // @[Cache_Soc.scala 89:22]
  reg  plru0_58; // @[Cache_Soc.scala 89:22]
  reg  plru0_59; // @[Cache_Soc.scala 89:22]
  reg  plru0_60; // @[Cache_Soc.scala 89:22]
  reg  plru0_61; // @[Cache_Soc.scala 89:22]
  reg  plru0_62; // @[Cache_Soc.scala 89:22]
  reg  plru0_63; // @[Cache_Soc.scala 89:22]
  reg  plru1_0; // @[Cache_Soc.scala 90:22]
  reg  plru1_1; // @[Cache_Soc.scala 90:22]
  reg  plru1_2; // @[Cache_Soc.scala 90:22]
  reg  plru1_3; // @[Cache_Soc.scala 90:22]
  reg  plru1_4; // @[Cache_Soc.scala 90:22]
  reg  plru1_5; // @[Cache_Soc.scala 90:22]
  reg  plru1_6; // @[Cache_Soc.scala 90:22]
  reg  plru1_7; // @[Cache_Soc.scala 90:22]
  reg  plru1_8; // @[Cache_Soc.scala 90:22]
  reg  plru1_9; // @[Cache_Soc.scala 90:22]
  reg  plru1_10; // @[Cache_Soc.scala 90:22]
  reg  plru1_11; // @[Cache_Soc.scala 90:22]
  reg  plru1_12; // @[Cache_Soc.scala 90:22]
  reg  plru1_13; // @[Cache_Soc.scala 90:22]
  reg  plru1_14; // @[Cache_Soc.scala 90:22]
  reg  plru1_15; // @[Cache_Soc.scala 90:22]
  reg  plru1_16; // @[Cache_Soc.scala 90:22]
  reg  plru1_17; // @[Cache_Soc.scala 90:22]
  reg  plru1_18; // @[Cache_Soc.scala 90:22]
  reg  plru1_19; // @[Cache_Soc.scala 90:22]
  reg  plru1_20; // @[Cache_Soc.scala 90:22]
  reg  plru1_21; // @[Cache_Soc.scala 90:22]
  reg  plru1_22; // @[Cache_Soc.scala 90:22]
  reg  plru1_23; // @[Cache_Soc.scala 90:22]
  reg  plru1_24; // @[Cache_Soc.scala 90:22]
  reg  plru1_25; // @[Cache_Soc.scala 90:22]
  reg  plru1_26; // @[Cache_Soc.scala 90:22]
  reg  plru1_27; // @[Cache_Soc.scala 90:22]
  reg  plru1_28; // @[Cache_Soc.scala 90:22]
  reg  plru1_29; // @[Cache_Soc.scala 90:22]
  reg  plru1_30; // @[Cache_Soc.scala 90:22]
  reg  plru1_31; // @[Cache_Soc.scala 90:22]
  reg  plru1_32; // @[Cache_Soc.scala 90:22]
  reg  plru1_33; // @[Cache_Soc.scala 90:22]
  reg  plru1_34; // @[Cache_Soc.scala 90:22]
  reg  plru1_35; // @[Cache_Soc.scala 90:22]
  reg  plru1_36; // @[Cache_Soc.scala 90:22]
  reg  plru1_37; // @[Cache_Soc.scala 90:22]
  reg  plru1_38; // @[Cache_Soc.scala 90:22]
  reg  plru1_39; // @[Cache_Soc.scala 90:22]
  reg  plru1_40; // @[Cache_Soc.scala 90:22]
  reg  plru1_41; // @[Cache_Soc.scala 90:22]
  reg  plru1_42; // @[Cache_Soc.scala 90:22]
  reg  plru1_43; // @[Cache_Soc.scala 90:22]
  reg  plru1_44; // @[Cache_Soc.scala 90:22]
  reg  plru1_45; // @[Cache_Soc.scala 90:22]
  reg  plru1_46; // @[Cache_Soc.scala 90:22]
  reg  plru1_47; // @[Cache_Soc.scala 90:22]
  reg  plru1_48; // @[Cache_Soc.scala 90:22]
  reg  plru1_49; // @[Cache_Soc.scala 90:22]
  reg  plru1_50; // @[Cache_Soc.scala 90:22]
  reg  plru1_51; // @[Cache_Soc.scala 90:22]
  reg  plru1_52; // @[Cache_Soc.scala 90:22]
  reg  plru1_53; // @[Cache_Soc.scala 90:22]
  reg  plru1_54; // @[Cache_Soc.scala 90:22]
  reg  plru1_55; // @[Cache_Soc.scala 90:22]
  reg  plru1_56; // @[Cache_Soc.scala 90:22]
  reg  plru1_57; // @[Cache_Soc.scala 90:22]
  reg  plru1_58; // @[Cache_Soc.scala 90:22]
  reg  plru1_59; // @[Cache_Soc.scala 90:22]
  reg  plru1_60; // @[Cache_Soc.scala 90:22]
  reg  plru1_61; // @[Cache_Soc.scala 90:22]
  reg  plru1_62; // @[Cache_Soc.scala 90:22]
  reg  plru1_63; // @[Cache_Soc.scala 90:22]
  reg  plru2_0; // @[Cache_Soc.scala 91:22]
  reg  plru2_1; // @[Cache_Soc.scala 91:22]
  reg  plru2_2; // @[Cache_Soc.scala 91:22]
  reg  plru2_3; // @[Cache_Soc.scala 91:22]
  reg  plru2_4; // @[Cache_Soc.scala 91:22]
  reg  plru2_5; // @[Cache_Soc.scala 91:22]
  reg  plru2_6; // @[Cache_Soc.scala 91:22]
  reg  plru2_7; // @[Cache_Soc.scala 91:22]
  reg  plru2_8; // @[Cache_Soc.scala 91:22]
  reg  plru2_9; // @[Cache_Soc.scala 91:22]
  reg  plru2_10; // @[Cache_Soc.scala 91:22]
  reg  plru2_11; // @[Cache_Soc.scala 91:22]
  reg  plru2_12; // @[Cache_Soc.scala 91:22]
  reg  plru2_13; // @[Cache_Soc.scala 91:22]
  reg  plru2_14; // @[Cache_Soc.scala 91:22]
  reg  plru2_15; // @[Cache_Soc.scala 91:22]
  reg  plru2_16; // @[Cache_Soc.scala 91:22]
  reg  plru2_17; // @[Cache_Soc.scala 91:22]
  reg  plru2_18; // @[Cache_Soc.scala 91:22]
  reg  plru2_19; // @[Cache_Soc.scala 91:22]
  reg  plru2_20; // @[Cache_Soc.scala 91:22]
  reg  plru2_21; // @[Cache_Soc.scala 91:22]
  reg  plru2_22; // @[Cache_Soc.scala 91:22]
  reg  plru2_23; // @[Cache_Soc.scala 91:22]
  reg  plru2_24; // @[Cache_Soc.scala 91:22]
  reg  plru2_25; // @[Cache_Soc.scala 91:22]
  reg  plru2_26; // @[Cache_Soc.scala 91:22]
  reg  plru2_27; // @[Cache_Soc.scala 91:22]
  reg  plru2_28; // @[Cache_Soc.scala 91:22]
  reg  plru2_29; // @[Cache_Soc.scala 91:22]
  reg  plru2_30; // @[Cache_Soc.scala 91:22]
  reg  plru2_31; // @[Cache_Soc.scala 91:22]
  reg  plru2_32; // @[Cache_Soc.scala 91:22]
  reg  plru2_33; // @[Cache_Soc.scala 91:22]
  reg  plru2_34; // @[Cache_Soc.scala 91:22]
  reg  plru2_35; // @[Cache_Soc.scala 91:22]
  reg  plru2_36; // @[Cache_Soc.scala 91:22]
  reg  plru2_37; // @[Cache_Soc.scala 91:22]
  reg  plru2_38; // @[Cache_Soc.scala 91:22]
  reg  plru2_39; // @[Cache_Soc.scala 91:22]
  reg  plru2_40; // @[Cache_Soc.scala 91:22]
  reg  plru2_41; // @[Cache_Soc.scala 91:22]
  reg  plru2_42; // @[Cache_Soc.scala 91:22]
  reg  plru2_43; // @[Cache_Soc.scala 91:22]
  reg  plru2_44; // @[Cache_Soc.scala 91:22]
  reg  plru2_45; // @[Cache_Soc.scala 91:22]
  reg  plru2_46; // @[Cache_Soc.scala 91:22]
  reg  plru2_47; // @[Cache_Soc.scala 91:22]
  reg  plru2_48; // @[Cache_Soc.scala 91:22]
  reg  plru2_49; // @[Cache_Soc.scala 91:22]
  reg  plru2_50; // @[Cache_Soc.scala 91:22]
  reg  plru2_51; // @[Cache_Soc.scala 91:22]
  reg  plru2_52; // @[Cache_Soc.scala 91:22]
  reg  plru2_53; // @[Cache_Soc.scala 91:22]
  reg  plru2_54; // @[Cache_Soc.scala 91:22]
  reg  plru2_55; // @[Cache_Soc.scala 91:22]
  reg  plru2_56; // @[Cache_Soc.scala 91:22]
  reg  plru2_57; // @[Cache_Soc.scala 91:22]
  reg  plru2_58; // @[Cache_Soc.scala 91:22]
  reg  plru2_59; // @[Cache_Soc.scala 91:22]
  reg  plru2_60; // @[Cache_Soc.scala 91:22]
  reg  plru2_61; // @[Cache_Soc.scala 91:22]
  reg  plru2_62; // @[Cache_Soc.scala 91:22]
  reg  plru2_63; // @[Cache_Soc.scala 91:22]
  wire  _T = state == 3'h1; // @[Cache_Soc.scala 94:16]
  wire  _T_1 = state == 3'h1 & cache_hit; // @[Cache_Soc.scala 94:28]
  wire  _GEN_0 = 6'h0 == rb_index ? hit_0 | hit_1 : plru0_0; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_1 = 6'h1 == rb_index ? hit_0 | hit_1 : plru0_1; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_2 = 6'h2 == rb_index ? hit_0 | hit_1 : plru0_2; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_3 = 6'h3 == rb_index ? hit_0 | hit_1 : plru0_3; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_4 = 6'h4 == rb_index ? hit_0 | hit_1 : plru0_4; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_5 = 6'h5 == rb_index ? hit_0 | hit_1 : plru0_5; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_6 = 6'h6 == rb_index ? hit_0 | hit_1 : plru0_6; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_7 = 6'h7 == rb_index ? hit_0 | hit_1 : plru0_7; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_8 = 6'h8 == rb_index ? hit_0 | hit_1 : plru0_8; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_9 = 6'h9 == rb_index ? hit_0 | hit_1 : plru0_9; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_10 = 6'ha == rb_index ? hit_0 | hit_1 : plru0_10; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_11 = 6'hb == rb_index ? hit_0 | hit_1 : plru0_11; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_12 = 6'hc == rb_index ? hit_0 | hit_1 : plru0_12; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_13 = 6'hd == rb_index ? hit_0 | hit_1 : plru0_13; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_14 = 6'he == rb_index ? hit_0 | hit_1 : plru0_14; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_15 = 6'hf == rb_index ? hit_0 | hit_1 : plru0_15; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_16 = 6'h10 == rb_index ? hit_0 | hit_1 : plru0_16; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_17 = 6'h11 == rb_index ? hit_0 | hit_1 : plru0_17; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_18 = 6'h12 == rb_index ? hit_0 | hit_1 : plru0_18; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_19 = 6'h13 == rb_index ? hit_0 | hit_1 : plru0_19; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_20 = 6'h14 == rb_index ? hit_0 | hit_1 : plru0_20; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_21 = 6'h15 == rb_index ? hit_0 | hit_1 : plru0_21; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_22 = 6'h16 == rb_index ? hit_0 | hit_1 : plru0_22; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_23 = 6'h17 == rb_index ? hit_0 | hit_1 : plru0_23; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_24 = 6'h18 == rb_index ? hit_0 | hit_1 : plru0_24; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_25 = 6'h19 == rb_index ? hit_0 | hit_1 : plru0_25; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_26 = 6'h1a == rb_index ? hit_0 | hit_1 : plru0_26; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_27 = 6'h1b == rb_index ? hit_0 | hit_1 : plru0_27; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_28 = 6'h1c == rb_index ? hit_0 | hit_1 : plru0_28; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_29 = 6'h1d == rb_index ? hit_0 | hit_1 : plru0_29; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_30 = 6'h1e == rb_index ? hit_0 | hit_1 : plru0_30; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_31 = 6'h1f == rb_index ? hit_0 | hit_1 : plru0_31; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_32 = 6'h20 == rb_index ? hit_0 | hit_1 : plru0_32; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_33 = 6'h21 == rb_index ? hit_0 | hit_1 : plru0_33; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_34 = 6'h22 == rb_index ? hit_0 | hit_1 : plru0_34; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_35 = 6'h23 == rb_index ? hit_0 | hit_1 : plru0_35; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_36 = 6'h24 == rb_index ? hit_0 | hit_1 : plru0_36; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_37 = 6'h25 == rb_index ? hit_0 | hit_1 : plru0_37; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_38 = 6'h26 == rb_index ? hit_0 | hit_1 : plru0_38; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_39 = 6'h27 == rb_index ? hit_0 | hit_1 : plru0_39; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_40 = 6'h28 == rb_index ? hit_0 | hit_1 : plru0_40; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_41 = 6'h29 == rb_index ? hit_0 | hit_1 : plru0_41; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_42 = 6'h2a == rb_index ? hit_0 | hit_1 : plru0_42; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_43 = 6'h2b == rb_index ? hit_0 | hit_1 : plru0_43; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_44 = 6'h2c == rb_index ? hit_0 | hit_1 : plru0_44; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_45 = 6'h2d == rb_index ? hit_0 | hit_1 : plru0_45; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_46 = 6'h2e == rb_index ? hit_0 | hit_1 : plru0_46; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_47 = 6'h2f == rb_index ? hit_0 | hit_1 : plru0_47; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_48 = 6'h30 == rb_index ? hit_0 | hit_1 : plru0_48; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_49 = 6'h31 == rb_index ? hit_0 | hit_1 : plru0_49; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_50 = 6'h32 == rb_index ? hit_0 | hit_1 : plru0_50; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_51 = 6'h33 == rb_index ? hit_0 | hit_1 : plru0_51; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_52 = 6'h34 == rb_index ? hit_0 | hit_1 : plru0_52; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_53 = 6'h35 == rb_index ? hit_0 | hit_1 : plru0_53; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_54 = 6'h36 == rb_index ? hit_0 | hit_1 : plru0_54; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_55 = 6'h37 == rb_index ? hit_0 | hit_1 : plru0_55; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_56 = 6'h38 == rb_index ? hit_0 | hit_1 : plru0_56; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_57 = 6'h39 == rb_index ? hit_0 | hit_1 : plru0_57; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_58 = 6'h3a == rb_index ? hit_0 | hit_1 : plru0_58; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_59 = 6'h3b == rb_index ? hit_0 | hit_1 : plru0_59; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_60 = 6'h3c == rb_index ? hit_0 | hit_1 : plru0_60; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_61 = 6'h3d == rb_index ? hit_0 | hit_1 : plru0_61; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_62 = 6'h3e == rb_index ? hit_0 | hit_1 : plru0_62; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_63 = 6'h3f == rb_index ? hit_0 | hit_1 : plru0_63; // @[Cache_Soc.scala 95:21 Cache_Soc.scala 95:21 Cache_Soc.scala 89:22]
  wire  _GEN_2439 = 6'h0 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_64 = 6'h0 == rb_index | plru1_0; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2440 = 6'h1 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_65 = 6'h1 == rb_index | plru1_1; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2441 = 6'h2 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_66 = 6'h2 == rb_index | plru1_2; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2442 = 6'h3 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_67 = 6'h3 == rb_index | plru1_3; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2443 = 6'h4 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_68 = 6'h4 == rb_index | plru1_4; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2444 = 6'h5 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_69 = 6'h5 == rb_index | plru1_5; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2445 = 6'h6 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_70 = 6'h6 == rb_index | plru1_6; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2446 = 6'h7 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_71 = 6'h7 == rb_index | plru1_7; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2447 = 6'h8 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_72 = 6'h8 == rb_index | plru1_8; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2448 = 6'h9 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_73 = 6'h9 == rb_index | plru1_9; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2449 = 6'ha == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_74 = 6'ha == rb_index | plru1_10; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2450 = 6'hb == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_75 = 6'hb == rb_index | plru1_11; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2451 = 6'hc == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_76 = 6'hc == rb_index | plru1_12; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2452 = 6'hd == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_77 = 6'hd == rb_index | plru1_13; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2453 = 6'he == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_78 = 6'he == rb_index | plru1_14; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2454 = 6'hf == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_79 = 6'hf == rb_index | plru1_15; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2455 = 6'h10 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_80 = 6'h10 == rb_index | plru1_16; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2456 = 6'h11 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_81 = 6'h11 == rb_index | plru1_17; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2457 = 6'h12 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_82 = 6'h12 == rb_index | plru1_18; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2458 = 6'h13 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_83 = 6'h13 == rb_index | plru1_19; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2459 = 6'h14 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_84 = 6'h14 == rb_index | plru1_20; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2460 = 6'h15 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_85 = 6'h15 == rb_index | plru1_21; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2461 = 6'h16 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_86 = 6'h16 == rb_index | plru1_22; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2462 = 6'h17 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_87 = 6'h17 == rb_index | plru1_23; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2463 = 6'h18 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_88 = 6'h18 == rb_index | plru1_24; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2464 = 6'h19 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_89 = 6'h19 == rb_index | plru1_25; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2465 = 6'h1a == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_90 = 6'h1a == rb_index | plru1_26; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2466 = 6'h1b == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_91 = 6'h1b == rb_index | plru1_27; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2467 = 6'h1c == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_92 = 6'h1c == rb_index | plru1_28; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2468 = 6'h1d == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_93 = 6'h1d == rb_index | plru1_29; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2469 = 6'h1e == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_94 = 6'h1e == rb_index | plru1_30; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2470 = 6'h1f == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_95 = 6'h1f == rb_index | plru1_31; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2471 = 6'h20 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_96 = 6'h20 == rb_index | plru1_32; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2472 = 6'h21 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_97 = 6'h21 == rb_index | plru1_33; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2473 = 6'h22 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_98 = 6'h22 == rb_index | plru1_34; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2474 = 6'h23 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_99 = 6'h23 == rb_index | plru1_35; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2475 = 6'h24 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_100 = 6'h24 == rb_index | plru1_36; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2476 = 6'h25 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_101 = 6'h25 == rb_index | plru1_37; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2477 = 6'h26 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_102 = 6'h26 == rb_index | plru1_38; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2478 = 6'h27 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_103 = 6'h27 == rb_index | plru1_39; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2479 = 6'h28 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_104 = 6'h28 == rb_index | plru1_40; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2480 = 6'h29 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_105 = 6'h29 == rb_index | plru1_41; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2481 = 6'h2a == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_106 = 6'h2a == rb_index | plru1_42; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2482 = 6'h2b == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_107 = 6'h2b == rb_index | plru1_43; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2483 = 6'h2c == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_108 = 6'h2c == rb_index | plru1_44; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2484 = 6'h2d == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_109 = 6'h2d == rb_index | plru1_45; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2485 = 6'h2e == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_110 = 6'h2e == rb_index | plru1_46; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2486 = 6'h2f == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_111 = 6'h2f == rb_index | plru1_47; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2487 = 6'h30 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_112 = 6'h30 == rb_index | plru1_48; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2488 = 6'h31 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_113 = 6'h31 == rb_index | plru1_49; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2489 = 6'h32 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_114 = 6'h32 == rb_index | plru1_50; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2490 = 6'h33 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_115 = 6'h33 == rb_index | plru1_51; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2491 = 6'h34 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_116 = 6'h34 == rb_index | plru1_52; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2492 = 6'h35 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_117 = 6'h35 == rb_index | plru1_53; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2493 = 6'h36 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_118 = 6'h36 == rb_index | plru1_54; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2494 = 6'h37 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_119 = 6'h37 == rb_index | plru1_55; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2495 = 6'h38 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_120 = 6'h38 == rb_index | plru1_56; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2496 = 6'h39 == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_121 = 6'h39 == rb_index | plru1_57; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2497 = 6'h3a == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_122 = 6'h3a == rb_index | plru1_58; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2498 = 6'h3b == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_123 = 6'h3b == rb_index | plru1_59; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2499 = 6'h3c == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_124 = 6'h3c == rb_index | plru1_60; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2500 = 6'h3d == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_125 = 6'h3d == rb_index | plru1_61; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2501 = 6'h3e == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_126 = 6'h3e == rb_index | plru1_62; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_2502 = 6'h3f == rb_index; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_127 = 6'h3f == rb_index | plru1_63; // @[Cache_Soc.scala 97:23 Cache_Soc.scala 97:23 Cache_Soc.scala 90:22]
  wire  _GEN_128 = 6'h0 == rb_index ? 1'h0 : plru1_0; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_129 = 6'h1 == rb_index ? 1'h0 : plru1_1; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_130 = 6'h2 == rb_index ? 1'h0 : plru1_2; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_131 = 6'h3 == rb_index ? 1'h0 : plru1_3; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_132 = 6'h4 == rb_index ? 1'h0 : plru1_4; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_133 = 6'h5 == rb_index ? 1'h0 : plru1_5; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_134 = 6'h6 == rb_index ? 1'h0 : plru1_6; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_135 = 6'h7 == rb_index ? 1'h0 : plru1_7; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_136 = 6'h8 == rb_index ? 1'h0 : plru1_8; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_137 = 6'h9 == rb_index ? 1'h0 : plru1_9; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_138 = 6'ha == rb_index ? 1'h0 : plru1_10; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_139 = 6'hb == rb_index ? 1'h0 : plru1_11; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_140 = 6'hc == rb_index ? 1'h0 : plru1_12; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_141 = 6'hd == rb_index ? 1'h0 : plru1_13; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_142 = 6'he == rb_index ? 1'h0 : plru1_14; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_143 = 6'hf == rb_index ? 1'h0 : plru1_15; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_144 = 6'h10 == rb_index ? 1'h0 : plru1_16; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_145 = 6'h11 == rb_index ? 1'h0 : plru1_17; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_146 = 6'h12 == rb_index ? 1'h0 : plru1_18; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_147 = 6'h13 == rb_index ? 1'h0 : plru1_19; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_148 = 6'h14 == rb_index ? 1'h0 : plru1_20; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_149 = 6'h15 == rb_index ? 1'h0 : plru1_21; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_150 = 6'h16 == rb_index ? 1'h0 : plru1_22; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_151 = 6'h17 == rb_index ? 1'h0 : plru1_23; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_152 = 6'h18 == rb_index ? 1'h0 : plru1_24; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_153 = 6'h19 == rb_index ? 1'h0 : plru1_25; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_154 = 6'h1a == rb_index ? 1'h0 : plru1_26; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_155 = 6'h1b == rb_index ? 1'h0 : plru1_27; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_156 = 6'h1c == rb_index ? 1'h0 : plru1_28; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_157 = 6'h1d == rb_index ? 1'h0 : plru1_29; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_158 = 6'h1e == rb_index ? 1'h0 : plru1_30; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_159 = 6'h1f == rb_index ? 1'h0 : plru1_31; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_160 = 6'h20 == rb_index ? 1'h0 : plru1_32; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_161 = 6'h21 == rb_index ? 1'h0 : plru1_33; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_162 = 6'h22 == rb_index ? 1'h0 : plru1_34; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_163 = 6'h23 == rb_index ? 1'h0 : plru1_35; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_164 = 6'h24 == rb_index ? 1'h0 : plru1_36; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_165 = 6'h25 == rb_index ? 1'h0 : plru1_37; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_166 = 6'h26 == rb_index ? 1'h0 : plru1_38; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_167 = 6'h27 == rb_index ? 1'h0 : plru1_39; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_168 = 6'h28 == rb_index ? 1'h0 : plru1_40; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_169 = 6'h29 == rb_index ? 1'h0 : plru1_41; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_170 = 6'h2a == rb_index ? 1'h0 : plru1_42; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_171 = 6'h2b == rb_index ? 1'h0 : plru1_43; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_172 = 6'h2c == rb_index ? 1'h0 : plru1_44; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_173 = 6'h2d == rb_index ? 1'h0 : plru1_45; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_174 = 6'h2e == rb_index ? 1'h0 : plru1_46; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_175 = 6'h2f == rb_index ? 1'h0 : plru1_47; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_176 = 6'h30 == rb_index ? 1'h0 : plru1_48; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_177 = 6'h31 == rb_index ? 1'h0 : plru1_49; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_178 = 6'h32 == rb_index ? 1'h0 : plru1_50; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_179 = 6'h33 == rb_index ? 1'h0 : plru1_51; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_180 = 6'h34 == rb_index ? 1'h0 : plru1_52; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_181 = 6'h35 == rb_index ? 1'h0 : plru1_53; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_182 = 6'h36 == rb_index ? 1'h0 : plru1_54; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_183 = 6'h37 == rb_index ? 1'h0 : plru1_55; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_184 = 6'h38 == rb_index ? 1'h0 : plru1_56; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_185 = 6'h39 == rb_index ? 1'h0 : plru1_57; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_186 = 6'h3a == rb_index ? 1'h0 : plru1_58; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_187 = 6'h3b == rb_index ? 1'h0 : plru1_59; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_188 = 6'h3c == rb_index ? 1'h0 : plru1_60; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_189 = 6'h3d == rb_index ? 1'h0 : plru1_61; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_190 = 6'h3e == rb_index ? 1'h0 : plru1_62; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_191 = 6'h3f == rb_index ? 1'h0 : plru1_63; // @[Cache_Soc.scala 99:23 Cache_Soc.scala 99:23 Cache_Soc.scala 90:22]
  wire  _GEN_192 = _GEN_2439 | plru2_0; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_193 = _GEN_2440 | plru2_1; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_194 = _GEN_2441 | plru2_2; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_195 = _GEN_2442 | plru2_3; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_196 = _GEN_2443 | plru2_4; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_197 = _GEN_2444 | plru2_5; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_198 = _GEN_2445 | plru2_6; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_199 = _GEN_2446 | plru2_7; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_200 = _GEN_2447 | plru2_8; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_201 = _GEN_2448 | plru2_9; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_202 = _GEN_2449 | plru2_10; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_203 = _GEN_2450 | plru2_11; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_204 = _GEN_2451 | plru2_12; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_205 = _GEN_2452 | plru2_13; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_206 = _GEN_2453 | plru2_14; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_207 = _GEN_2454 | plru2_15; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_208 = _GEN_2455 | plru2_16; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_209 = _GEN_2456 | plru2_17; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_210 = _GEN_2457 | plru2_18; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_211 = _GEN_2458 | plru2_19; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_212 = _GEN_2459 | plru2_20; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_213 = _GEN_2460 | plru2_21; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_214 = _GEN_2461 | plru2_22; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_215 = _GEN_2462 | plru2_23; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_216 = _GEN_2463 | plru2_24; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_217 = _GEN_2464 | plru2_25; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_218 = _GEN_2465 | plru2_26; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_219 = _GEN_2466 | plru2_27; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_220 = _GEN_2467 | plru2_28; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_221 = _GEN_2468 | plru2_29; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_222 = _GEN_2469 | plru2_30; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_223 = _GEN_2470 | plru2_31; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_224 = _GEN_2471 | plru2_32; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_225 = _GEN_2472 | plru2_33; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_226 = _GEN_2473 | plru2_34; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_227 = _GEN_2474 | plru2_35; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_228 = _GEN_2475 | plru2_36; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_229 = _GEN_2476 | plru2_37; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_230 = _GEN_2477 | plru2_38; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_231 = _GEN_2478 | plru2_39; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_232 = _GEN_2479 | plru2_40; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_233 = _GEN_2480 | plru2_41; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_234 = _GEN_2481 | plru2_42; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_235 = _GEN_2482 | plru2_43; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_236 = _GEN_2483 | plru2_44; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_237 = _GEN_2484 | plru2_45; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_238 = _GEN_2485 | plru2_46; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_239 = _GEN_2486 | plru2_47; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_240 = _GEN_2487 | plru2_48; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_241 = _GEN_2488 | plru2_49; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_242 = _GEN_2489 | plru2_50; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_243 = _GEN_2490 | plru2_51; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_244 = _GEN_2491 | plru2_52; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_245 = _GEN_2492 | plru2_53; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_246 = _GEN_2493 | plru2_54; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_247 = _GEN_2494 | plru2_55; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_248 = _GEN_2495 | plru2_56; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_249 = _GEN_2496 | plru2_57; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_250 = _GEN_2497 | plru2_58; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_251 = _GEN_2498 | plru2_59; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_252 = _GEN_2499 | plru2_60; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_253 = _GEN_2500 | plru2_61; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_254 = _GEN_2501 | plru2_62; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_255 = _GEN_2502 | plru2_63; // @[Cache_Soc.scala 101:23 Cache_Soc.scala 101:23 Cache_Soc.scala 91:22]
  wire  _GEN_256 = 6'h0 == rb_index ? 1'h0 : plru2_0; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_257 = 6'h1 == rb_index ? 1'h0 : plru2_1; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_258 = 6'h2 == rb_index ? 1'h0 : plru2_2; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_259 = 6'h3 == rb_index ? 1'h0 : plru2_3; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_260 = 6'h4 == rb_index ? 1'h0 : plru2_4; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_261 = 6'h5 == rb_index ? 1'h0 : plru2_5; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_262 = 6'h6 == rb_index ? 1'h0 : plru2_6; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_263 = 6'h7 == rb_index ? 1'h0 : plru2_7; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_264 = 6'h8 == rb_index ? 1'h0 : plru2_8; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_265 = 6'h9 == rb_index ? 1'h0 : plru2_9; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_266 = 6'ha == rb_index ? 1'h0 : plru2_10; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_267 = 6'hb == rb_index ? 1'h0 : plru2_11; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_268 = 6'hc == rb_index ? 1'h0 : plru2_12; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_269 = 6'hd == rb_index ? 1'h0 : plru2_13; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_270 = 6'he == rb_index ? 1'h0 : plru2_14; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_271 = 6'hf == rb_index ? 1'h0 : plru2_15; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_272 = 6'h10 == rb_index ? 1'h0 : plru2_16; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_273 = 6'h11 == rb_index ? 1'h0 : plru2_17; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_274 = 6'h12 == rb_index ? 1'h0 : plru2_18; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_275 = 6'h13 == rb_index ? 1'h0 : plru2_19; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_276 = 6'h14 == rb_index ? 1'h0 : plru2_20; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_277 = 6'h15 == rb_index ? 1'h0 : plru2_21; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_278 = 6'h16 == rb_index ? 1'h0 : plru2_22; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_279 = 6'h17 == rb_index ? 1'h0 : plru2_23; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_280 = 6'h18 == rb_index ? 1'h0 : plru2_24; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_281 = 6'h19 == rb_index ? 1'h0 : plru2_25; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_282 = 6'h1a == rb_index ? 1'h0 : plru2_26; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_283 = 6'h1b == rb_index ? 1'h0 : plru2_27; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_284 = 6'h1c == rb_index ? 1'h0 : plru2_28; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_285 = 6'h1d == rb_index ? 1'h0 : plru2_29; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_286 = 6'h1e == rb_index ? 1'h0 : plru2_30; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_287 = 6'h1f == rb_index ? 1'h0 : plru2_31; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_288 = 6'h20 == rb_index ? 1'h0 : plru2_32; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_289 = 6'h21 == rb_index ? 1'h0 : plru2_33; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_290 = 6'h22 == rb_index ? 1'h0 : plru2_34; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_291 = 6'h23 == rb_index ? 1'h0 : plru2_35; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_292 = 6'h24 == rb_index ? 1'h0 : plru2_36; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_293 = 6'h25 == rb_index ? 1'h0 : plru2_37; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_294 = 6'h26 == rb_index ? 1'h0 : plru2_38; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_295 = 6'h27 == rb_index ? 1'h0 : plru2_39; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_296 = 6'h28 == rb_index ? 1'h0 : plru2_40; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_297 = 6'h29 == rb_index ? 1'h0 : plru2_41; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_298 = 6'h2a == rb_index ? 1'h0 : plru2_42; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_299 = 6'h2b == rb_index ? 1'h0 : plru2_43; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_300 = 6'h2c == rb_index ? 1'h0 : plru2_44; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_301 = 6'h2d == rb_index ? 1'h0 : plru2_45; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_302 = 6'h2e == rb_index ? 1'h0 : plru2_46; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_303 = 6'h2f == rb_index ? 1'h0 : plru2_47; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_304 = 6'h30 == rb_index ? 1'h0 : plru2_48; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_305 = 6'h31 == rb_index ? 1'h0 : plru2_49; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_306 = 6'h32 == rb_index ? 1'h0 : plru2_50; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_307 = 6'h33 == rb_index ? 1'h0 : plru2_51; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_308 = 6'h34 == rb_index ? 1'h0 : plru2_52; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_309 = 6'h35 == rb_index ? 1'h0 : plru2_53; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_310 = 6'h36 == rb_index ? 1'h0 : plru2_54; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_311 = 6'h37 == rb_index ? 1'h0 : plru2_55; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_312 = 6'h38 == rb_index ? 1'h0 : plru2_56; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_313 = 6'h39 == rb_index ? 1'h0 : plru2_57; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_314 = 6'h3a == rb_index ? 1'h0 : plru2_58; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_315 = 6'h3b == rb_index ? 1'h0 : plru2_59; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_316 = 6'h3c == rb_index ? 1'h0 : plru2_60; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_317 = 6'h3d == rb_index ? 1'h0 : plru2_61; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_318 = 6'h3e == rb_index ? 1'h0 : plru2_62; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_319 = 6'h3f == rb_index ? 1'h0 : plru2_63; // @[Cache_Soc.scala 103:23 Cache_Soc.scala 103:23 Cache_Soc.scala 91:22]
  wire  _GEN_320 = hit_3 ? _GEN_256 : plru2_0; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_321 = hit_3 ? _GEN_257 : plru2_1; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_322 = hit_3 ? _GEN_258 : plru2_2; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_323 = hit_3 ? _GEN_259 : plru2_3; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_324 = hit_3 ? _GEN_260 : plru2_4; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_325 = hit_3 ? _GEN_261 : plru2_5; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_326 = hit_3 ? _GEN_262 : plru2_6; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_327 = hit_3 ? _GEN_263 : plru2_7; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_328 = hit_3 ? _GEN_264 : plru2_8; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_329 = hit_3 ? _GEN_265 : plru2_9; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_330 = hit_3 ? _GEN_266 : plru2_10; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_331 = hit_3 ? _GEN_267 : plru2_11; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_332 = hit_3 ? _GEN_268 : plru2_12; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_333 = hit_3 ? _GEN_269 : plru2_13; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_334 = hit_3 ? _GEN_270 : plru2_14; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_335 = hit_3 ? _GEN_271 : plru2_15; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_336 = hit_3 ? _GEN_272 : plru2_16; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_337 = hit_3 ? _GEN_273 : plru2_17; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_338 = hit_3 ? _GEN_274 : plru2_18; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_339 = hit_3 ? _GEN_275 : plru2_19; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_340 = hit_3 ? _GEN_276 : plru2_20; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_341 = hit_3 ? _GEN_277 : plru2_21; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_342 = hit_3 ? _GEN_278 : plru2_22; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_343 = hit_3 ? _GEN_279 : plru2_23; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_344 = hit_3 ? _GEN_280 : plru2_24; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_345 = hit_3 ? _GEN_281 : plru2_25; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_346 = hit_3 ? _GEN_282 : plru2_26; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_347 = hit_3 ? _GEN_283 : plru2_27; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_348 = hit_3 ? _GEN_284 : plru2_28; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_349 = hit_3 ? _GEN_285 : plru2_29; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_350 = hit_3 ? _GEN_286 : plru2_30; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_351 = hit_3 ? _GEN_287 : plru2_31; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_352 = hit_3 ? _GEN_288 : plru2_32; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_353 = hit_3 ? _GEN_289 : plru2_33; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_354 = hit_3 ? _GEN_290 : plru2_34; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_355 = hit_3 ? _GEN_291 : plru2_35; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_356 = hit_3 ? _GEN_292 : plru2_36; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_357 = hit_3 ? _GEN_293 : plru2_37; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_358 = hit_3 ? _GEN_294 : plru2_38; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_359 = hit_3 ? _GEN_295 : plru2_39; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_360 = hit_3 ? _GEN_296 : plru2_40; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_361 = hit_3 ? _GEN_297 : plru2_41; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_362 = hit_3 ? _GEN_298 : plru2_42; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_363 = hit_3 ? _GEN_299 : plru2_43; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_364 = hit_3 ? _GEN_300 : plru2_44; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_365 = hit_3 ? _GEN_301 : plru2_45; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_366 = hit_3 ? _GEN_302 : plru2_46; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_367 = hit_3 ? _GEN_303 : plru2_47; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_368 = hit_3 ? _GEN_304 : plru2_48; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_369 = hit_3 ? _GEN_305 : plru2_49; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_370 = hit_3 ? _GEN_306 : plru2_50; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_371 = hit_3 ? _GEN_307 : plru2_51; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_372 = hit_3 ? _GEN_308 : plru2_52; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_373 = hit_3 ? _GEN_309 : plru2_53; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_374 = hit_3 ? _GEN_310 : plru2_54; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_375 = hit_3 ? _GEN_311 : plru2_55; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_376 = hit_3 ? _GEN_312 : plru2_56; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_377 = hit_3 ? _GEN_313 : plru2_57; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_378 = hit_3 ? _GEN_314 : plru2_58; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_379 = hit_3 ? _GEN_315 : plru2_59; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_380 = hit_3 ? _GEN_316 : plru2_60; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_381 = hit_3 ? _GEN_317 : plru2_61; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_382 = hit_3 ? _GEN_318 : plru2_62; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_383 = hit_3 ? _GEN_319 : plru2_63; // @[Cache_Soc.scala 102:26 Cache_Soc.scala 91:22]
  wire  _GEN_384 = hit_2 ? _GEN_192 : _GEN_320; // @[Cache_Soc.scala 100:26]
  wire  _GEN_385 = hit_2 ? _GEN_193 : _GEN_321; // @[Cache_Soc.scala 100:26]
  wire  _GEN_386 = hit_2 ? _GEN_194 : _GEN_322; // @[Cache_Soc.scala 100:26]
  wire  _GEN_387 = hit_2 ? _GEN_195 : _GEN_323; // @[Cache_Soc.scala 100:26]
  wire  _GEN_388 = hit_2 ? _GEN_196 : _GEN_324; // @[Cache_Soc.scala 100:26]
  wire  _GEN_389 = hit_2 ? _GEN_197 : _GEN_325; // @[Cache_Soc.scala 100:26]
  wire  _GEN_390 = hit_2 ? _GEN_198 : _GEN_326; // @[Cache_Soc.scala 100:26]
  wire  _GEN_391 = hit_2 ? _GEN_199 : _GEN_327; // @[Cache_Soc.scala 100:26]
  wire  _GEN_392 = hit_2 ? _GEN_200 : _GEN_328; // @[Cache_Soc.scala 100:26]
  wire  _GEN_393 = hit_2 ? _GEN_201 : _GEN_329; // @[Cache_Soc.scala 100:26]
  wire  _GEN_394 = hit_2 ? _GEN_202 : _GEN_330; // @[Cache_Soc.scala 100:26]
  wire  _GEN_395 = hit_2 ? _GEN_203 : _GEN_331; // @[Cache_Soc.scala 100:26]
  wire  _GEN_396 = hit_2 ? _GEN_204 : _GEN_332; // @[Cache_Soc.scala 100:26]
  wire  _GEN_397 = hit_2 ? _GEN_205 : _GEN_333; // @[Cache_Soc.scala 100:26]
  wire  _GEN_398 = hit_2 ? _GEN_206 : _GEN_334; // @[Cache_Soc.scala 100:26]
  wire  _GEN_399 = hit_2 ? _GEN_207 : _GEN_335; // @[Cache_Soc.scala 100:26]
  wire  _GEN_400 = hit_2 ? _GEN_208 : _GEN_336; // @[Cache_Soc.scala 100:26]
  wire  _GEN_401 = hit_2 ? _GEN_209 : _GEN_337; // @[Cache_Soc.scala 100:26]
  wire  _GEN_402 = hit_2 ? _GEN_210 : _GEN_338; // @[Cache_Soc.scala 100:26]
  wire  _GEN_403 = hit_2 ? _GEN_211 : _GEN_339; // @[Cache_Soc.scala 100:26]
  wire  _GEN_404 = hit_2 ? _GEN_212 : _GEN_340; // @[Cache_Soc.scala 100:26]
  wire  _GEN_405 = hit_2 ? _GEN_213 : _GEN_341; // @[Cache_Soc.scala 100:26]
  wire  _GEN_406 = hit_2 ? _GEN_214 : _GEN_342; // @[Cache_Soc.scala 100:26]
  wire  _GEN_407 = hit_2 ? _GEN_215 : _GEN_343; // @[Cache_Soc.scala 100:26]
  wire  _GEN_408 = hit_2 ? _GEN_216 : _GEN_344; // @[Cache_Soc.scala 100:26]
  wire  _GEN_409 = hit_2 ? _GEN_217 : _GEN_345; // @[Cache_Soc.scala 100:26]
  wire  _GEN_410 = hit_2 ? _GEN_218 : _GEN_346; // @[Cache_Soc.scala 100:26]
  wire  _GEN_411 = hit_2 ? _GEN_219 : _GEN_347; // @[Cache_Soc.scala 100:26]
  wire  _GEN_412 = hit_2 ? _GEN_220 : _GEN_348; // @[Cache_Soc.scala 100:26]
  wire  _GEN_413 = hit_2 ? _GEN_221 : _GEN_349; // @[Cache_Soc.scala 100:26]
  wire  _GEN_414 = hit_2 ? _GEN_222 : _GEN_350; // @[Cache_Soc.scala 100:26]
  wire  _GEN_415 = hit_2 ? _GEN_223 : _GEN_351; // @[Cache_Soc.scala 100:26]
  wire  _GEN_416 = hit_2 ? _GEN_224 : _GEN_352; // @[Cache_Soc.scala 100:26]
  wire  _GEN_417 = hit_2 ? _GEN_225 : _GEN_353; // @[Cache_Soc.scala 100:26]
  wire  _GEN_418 = hit_2 ? _GEN_226 : _GEN_354; // @[Cache_Soc.scala 100:26]
  wire  _GEN_419 = hit_2 ? _GEN_227 : _GEN_355; // @[Cache_Soc.scala 100:26]
  wire  _GEN_420 = hit_2 ? _GEN_228 : _GEN_356; // @[Cache_Soc.scala 100:26]
  wire  _GEN_421 = hit_2 ? _GEN_229 : _GEN_357; // @[Cache_Soc.scala 100:26]
  wire  _GEN_422 = hit_2 ? _GEN_230 : _GEN_358; // @[Cache_Soc.scala 100:26]
  wire  _GEN_423 = hit_2 ? _GEN_231 : _GEN_359; // @[Cache_Soc.scala 100:26]
  wire  _GEN_424 = hit_2 ? _GEN_232 : _GEN_360; // @[Cache_Soc.scala 100:26]
  wire  _GEN_425 = hit_2 ? _GEN_233 : _GEN_361; // @[Cache_Soc.scala 100:26]
  wire  _GEN_426 = hit_2 ? _GEN_234 : _GEN_362; // @[Cache_Soc.scala 100:26]
  wire  _GEN_427 = hit_2 ? _GEN_235 : _GEN_363; // @[Cache_Soc.scala 100:26]
  wire  _GEN_428 = hit_2 ? _GEN_236 : _GEN_364; // @[Cache_Soc.scala 100:26]
  wire  _GEN_429 = hit_2 ? _GEN_237 : _GEN_365; // @[Cache_Soc.scala 100:26]
  wire  _GEN_430 = hit_2 ? _GEN_238 : _GEN_366; // @[Cache_Soc.scala 100:26]
  wire  _GEN_431 = hit_2 ? _GEN_239 : _GEN_367; // @[Cache_Soc.scala 100:26]
  wire  _GEN_432 = hit_2 ? _GEN_240 : _GEN_368; // @[Cache_Soc.scala 100:26]
  wire  _GEN_433 = hit_2 ? _GEN_241 : _GEN_369; // @[Cache_Soc.scala 100:26]
  wire  _GEN_434 = hit_2 ? _GEN_242 : _GEN_370; // @[Cache_Soc.scala 100:26]
  wire  _GEN_435 = hit_2 ? _GEN_243 : _GEN_371; // @[Cache_Soc.scala 100:26]
  wire  _GEN_436 = hit_2 ? _GEN_244 : _GEN_372; // @[Cache_Soc.scala 100:26]
  wire  _GEN_437 = hit_2 ? _GEN_245 : _GEN_373; // @[Cache_Soc.scala 100:26]
  wire  _GEN_438 = hit_2 ? _GEN_246 : _GEN_374; // @[Cache_Soc.scala 100:26]
  wire  _GEN_439 = hit_2 ? _GEN_247 : _GEN_375; // @[Cache_Soc.scala 100:26]
  wire  _GEN_440 = hit_2 ? _GEN_248 : _GEN_376; // @[Cache_Soc.scala 100:26]
  wire  _GEN_441 = hit_2 ? _GEN_249 : _GEN_377; // @[Cache_Soc.scala 100:26]
  wire  _GEN_442 = hit_2 ? _GEN_250 : _GEN_378; // @[Cache_Soc.scala 100:26]
  wire  _GEN_443 = hit_2 ? _GEN_251 : _GEN_379; // @[Cache_Soc.scala 100:26]
  wire  _GEN_444 = hit_2 ? _GEN_252 : _GEN_380; // @[Cache_Soc.scala 100:26]
  wire  _GEN_445 = hit_2 ? _GEN_253 : _GEN_381; // @[Cache_Soc.scala 100:26]
  wire  _GEN_446 = hit_2 ? _GEN_254 : _GEN_382; // @[Cache_Soc.scala 100:26]
  wire  _GEN_447 = hit_2 ? _GEN_255 : _GEN_383; // @[Cache_Soc.scala 100:26]
  wire  _GEN_448 = hit_1 ? _GEN_128 : plru1_0; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_449 = hit_1 ? _GEN_129 : plru1_1; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_450 = hit_1 ? _GEN_130 : plru1_2; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_451 = hit_1 ? _GEN_131 : plru1_3; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_452 = hit_1 ? _GEN_132 : plru1_4; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_453 = hit_1 ? _GEN_133 : plru1_5; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_454 = hit_1 ? _GEN_134 : plru1_6; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_455 = hit_1 ? _GEN_135 : plru1_7; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_456 = hit_1 ? _GEN_136 : plru1_8; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_457 = hit_1 ? _GEN_137 : plru1_9; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_458 = hit_1 ? _GEN_138 : plru1_10; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_459 = hit_1 ? _GEN_139 : plru1_11; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_460 = hit_1 ? _GEN_140 : plru1_12; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_461 = hit_1 ? _GEN_141 : plru1_13; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_462 = hit_1 ? _GEN_142 : plru1_14; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_463 = hit_1 ? _GEN_143 : plru1_15; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_464 = hit_1 ? _GEN_144 : plru1_16; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_465 = hit_1 ? _GEN_145 : plru1_17; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_466 = hit_1 ? _GEN_146 : plru1_18; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_467 = hit_1 ? _GEN_147 : plru1_19; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_468 = hit_1 ? _GEN_148 : plru1_20; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_469 = hit_1 ? _GEN_149 : plru1_21; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_470 = hit_1 ? _GEN_150 : plru1_22; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_471 = hit_1 ? _GEN_151 : plru1_23; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_472 = hit_1 ? _GEN_152 : plru1_24; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_473 = hit_1 ? _GEN_153 : plru1_25; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_474 = hit_1 ? _GEN_154 : plru1_26; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_475 = hit_1 ? _GEN_155 : plru1_27; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_476 = hit_1 ? _GEN_156 : plru1_28; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_477 = hit_1 ? _GEN_157 : plru1_29; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_478 = hit_1 ? _GEN_158 : plru1_30; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_479 = hit_1 ? _GEN_159 : plru1_31; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_480 = hit_1 ? _GEN_160 : plru1_32; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_481 = hit_1 ? _GEN_161 : plru1_33; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_482 = hit_1 ? _GEN_162 : plru1_34; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_483 = hit_1 ? _GEN_163 : plru1_35; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_484 = hit_1 ? _GEN_164 : plru1_36; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_485 = hit_1 ? _GEN_165 : plru1_37; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_486 = hit_1 ? _GEN_166 : plru1_38; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_487 = hit_1 ? _GEN_167 : plru1_39; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_488 = hit_1 ? _GEN_168 : plru1_40; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_489 = hit_1 ? _GEN_169 : plru1_41; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_490 = hit_1 ? _GEN_170 : plru1_42; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_491 = hit_1 ? _GEN_171 : plru1_43; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_492 = hit_1 ? _GEN_172 : plru1_44; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_493 = hit_1 ? _GEN_173 : plru1_45; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_494 = hit_1 ? _GEN_174 : plru1_46; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_495 = hit_1 ? _GEN_175 : plru1_47; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_496 = hit_1 ? _GEN_176 : plru1_48; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_497 = hit_1 ? _GEN_177 : plru1_49; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_498 = hit_1 ? _GEN_178 : plru1_50; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_499 = hit_1 ? _GEN_179 : plru1_51; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_500 = hit_1 ? _GEN_180 : plru1_52; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_501 = hit_1 ? _GEN_181 : plru1_53; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_502 = hit_1 ? _GEN_182 : plru1_54; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_503 = hit_1 ? _GEN_183 : plru1_55; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_504 = hit_1 ? _GEN_184 : plru1_56; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_505 = hit_1 ? _GEN_185 : plru1_57; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_506 = hit_1 ? _GEN_186 : plru1_58; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_507 = hit_1 ? _GEN_187 : plru1_59; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_508 = hit_1 ? _GEN_188 : plru1_60; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_509 = hit_1 ? _GEN_189 : plru1_61; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_510 = hit_1 ? _GEN_190 : plru1_62; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_511 = hit_1 ? _GEN_191 : plru1_63; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 90:22]
  wire  _GEN_512 = hit_1 ? plru2_0 : _GEN_384; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_513 = hit_1 ? plru2_1 : _GEN_385; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_514 = hit_1 ? plru2_2 : _GEN_386; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_515 = hit_1 ? plru2_3 : _GEN_387; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_516 = hit_1 ? plru2_4 : _GEN_388; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_517 = hit_1 ? plru2_5 : _GEN_389; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_518 = hit_1 ? plru2_6 : _GEN_390; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_519 = hit_1 ? plru2_7 : _GEN_391; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_520 = hit_1 ? plru2_8 : _GEN_392; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_521 = hit_1 ? plru2_9 : _GEN_393; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_522 = hit_1 ? plru2_10 : _GEN_394; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_523 = hit_1 ? plru2_11 : _GEN_395; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_524 = hit_1 ? plru2_12 : _GEN_396; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_525 = hit_1 ? plru2_13 : _GEN_397; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_526 = hit_1 ? plru2_14 : _GEN_398; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_527 = hit_1 ? plru2_15 : _GEN_399; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_528 = hit_1 ? plru2_16 : _GEN_400; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_529 = hit_1 ? plru2_17 : _GEN_401; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_530 = hit_1 ? plru2_18 : _GEN_402; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_531 = hit_1 ? plru2_19 : _GEN_403; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_532 = hit_1 ? plru2_20 : _GEN_404; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_533 = hit_1 ? plru2_21 : _GEN_405; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_534 = hit_1 ? plru2_22 : _GEN_406; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_535 = hit_1 ? plru2_23 : _GEN_407; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_536 = hit_1 ? plru2_24 : _GEN_408; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_537 = hit_1 ? plru2_25 : _GEN_409; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_538 = hit_1 ? plru2_26 : _GEN_410; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_539 = hit_1 ? plru2_27 : _GEN_411; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_540 = hit_1 ? plru2_28 : _GEN_412; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_541 = hit_1 ? plru2_29 : _GEN_413; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_542 = hit_1 ? plru2_30 : _GEN_414; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_543 = hit_1 ? plru2_31 : _GEN_415; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_544 = hit_1 ? plru2_32 : _GEN_416; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_545 = hit_1 ? plru2_33 : _GEN_417; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_546 = hit_1 ? plru2_34 : _GEN_418; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_547 = hit_1 ? plru2_35 : _GEN_419; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_548 = hit_1 ? plru2_36 : _GEN_420; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_549 = hit_1 ? plru2_37 : _GEN_421; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_550 = hit_1 ? plru2_38 : _GEN_422; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_551 = hit_1 ? plru2_39 : _GEN_423; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_552 = hit_1 ? plru2_40 : _GEN_424; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_553 = hit_1 ? plru2_41 : _GEN_425; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_554 = hit_1 ? plru2_42 : _GEN_426; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_555 = hit_1 ? plru2_43 : _GEN_427; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_556 = hit_1 ? plru2_44 : _GEN_428; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_557 = hit_1 ? plru2_45 : _GEN_429; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_558 = hit_1 ? plru2_46 : _GEN_430; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_559 = hit_1 ? plru2_47 : _GEN_431; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_560 = hit_1 ? plru2_48 : _GEN_432; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_561 = hit_1 ? plru2_49 : _GEN_433; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_562 = hit_1 ? plru2_50 : _GEN_434; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_563 = hit_1 ? plru2_51 : _GEN_435; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_564 = hit_1 ? plru2_52 : _GEN_436; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_565 = hit_1 ? plru2_53 : _GEN_437; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_566 = hit_1 ? plru2_54 : _GEN_438; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_567 = hit_1 ? plru2_55 : _GEN_439; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_568 = hit_1 ? plru2_56 : _GEN_440; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_569 = hit_1 ? plru2_57 : _GEN_441; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_570 = hit_1 ? plru2_58 : _GEN_442; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_571 = hit_1 ? plru2_59 : _GEN_443; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_572 = hit_1 ? plru2_60 : _GEN_444; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_573 = hit_1 ? plru2_61 : _GEN_445; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_574 = hit_1 ? plru2_62 : _GEN_446; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_575 = hit_1 ? plru2_63 : _GEN_447; // @[Cache_Soc.scala 98:26 Cache_Soc.scala 91:22]
  wire  _GEN_576 = hit_0 ? _GEN_64 : _GEN_448; // @[Cache_Soc.scala 96:19]
  wire  _GEN_577 = hit_0 ? _GEN_65 : _GEN_449; // @[Cache_Soc.scala 96:19]
  wire  _GEN_578 = hit_0 ? _GEN_66 : _GEN_450; // @[Cache_Soc.scala 96:19]
  wire  _GEN_579 = hit_0 ? _GEN_67 : _GEN_451; // @[Cache_Soc.scala 96:19]
  wire  _GEN_580 = hit_0 ? _GEN_68 : _GEN_452; // @[Cache_Soc.scala 96:19]
  wire  _GEN_581 = hit_0 ? _GEN_69 : _GEN_453; // @[Cache_Soc.scala 96:19]
  wire  _GEN_582 = hit_0 ? _GEN_70 : _GEN_454; // @[Cache_Soc.scala 96:19]
  wire  _GEN_583 = hit_0 ? _GEN_71 : _GEN_455; // @[Cache_Soc.scala 96:19]
  wire  _GEN_584 = hit_0 ? _GEN_72 : _GEN_456; // @[Cache_Soc.scala 96:19]
  wire  _GEN_585 = hit_0 ? _GEN_73 : _GEN_457; // @[Cache_Soc.scala 96:19]
  wire  _GEN_586 = hit_0 ? _GEN_74 : _GEN_458; // @[Cache_Soc.scala 96:19]
  wire  _GEN_587 = hit_0 ? _GEN_75 : _GEN_459; // @[Cache_Soc.scala 96:19]
  wire  _GEN_588 = hit_0 ? _GEN_76 : _GEN_460; // @[Cache_Soc.scala 96:19]
  wire  _GEN_589 = hit_0 ? _GEN_77 : _GEN_461; // @[Cache_Soc.scala 96:19]
  wire  _GEN_590 = hit_0 ? _GEN_78 : _GEN_462; // @[Cache_Soc.scala 96:19]
  wire  _GEN_591 = hit_0 ? _GEN_79 : _GEN_463; // @[Cache_Soc.scala 96:19]
  wire  _GEN_592 = hit_0 ? _GEN_80 : _GEN_464; // @[Cache_Soc.scala 96:19]
  wire  _GEN_593 = hit_0 ? _GEN_81 : _GEN_465; // @[Cache_Soc.scala 96:19]
  wire  _GEN_594 = hit_0 ? _GEN_82 : _GEN_466; // @[Cache_Soc.scala 96:19]
  wire  _GEN_595 = hit_0 ? _GEN_83 : _GEN_467; // @[Cache_Soc.scala 96:19]
  wire  _GEN_596 = hit_0 ? _GEN_84 : _GEN_468; // @[Cache_Soc.scala 96:19]
  wire  _GEN_597 = hit_0 ? _GEN_85 : _GEN_469; // @[Cache_Soc.scala 96:19]
  wire  _GEN_598 = hit_0 ? _GEN_86 : _GEN_470; // @[Cache_Soc.scala 96:19]
  wire  _GEN_599 = hit_0 ? _GEN_87 : _GEN_471; // @[Cache_Soc.scala 96:19]
  wire  _GEN_600 = hit_0 ? _GEN_88 : _GEN_472; // @[Cache_Soc.scala 96:19]
  wire  _GEN_601 = hit_0 ? _GEN_89 : _GEN_473; // @[Cache_Soc.scala 96:19]
  wire  _GEN_602 = hit_0 ? _GEN_90 : _GEN_474; // @[Cache_Soc.scala 96:19]
  wire  _GEN_603 = hit_0 ? _GEN_91 : _GEN_475; // @[Cache_Soc.scala 96:19]
  wire  _GEN_604 = hit_0 ? _GEN_92 : _GEN_476; // @[Cache_Soc.scala 96:19]
  wire  _GEN_605 = hit_0 ? _GEN_93 : _GEN_477; // @[Cache_Soc.scala 96:19]
  wire  _GEN_606 = hit_0 ? _GEN_94 : _GEN_478; // @[Cache_Soc.scala 96:19]
  wire  _GEN_607 = hit_0 ? _GEN_95 : _GEN_479; // @[Cache_Soc.scala 96:19]
  wire  _GEN_608 = hit_0 ? _GEN_96 : _GEN_480; // @[Cache_Soc.scala 96:19]
  wire  _GEN_609 = hit_0 ? _GEN_97 : _GEN_481; // @[Cache_Soc.scala 96:19]
  wire  _GEN_610 = hit_0 ? _GEN_98 : _GEN_482; // @[Cache_Soc.scala 96:19]
  wire  _GEN_611 = hit_0 ? _GEN_99 : _GEN_483; // @[Cache_Soc.scala 96:19]
  wire  _GEN_612 = hit_0 ? _GEN_100 : _GEN_484; // @[Cache_Soc.scala 96:19]
  wire  _GEN_613 = hit_0 ? _GEN_101 : _GEN_485; // @[Cache_Soc.scala 96:19]
  wire  _GEN_614 = hit_0 ? _GEN_102 : _GEN_486; // @[Cache_Soc.scala 96:19]
  wire  _GEN_615 = hit_0 ? _GEN_103 : _GEN_487; // @[Cache_Soc.scala 96:19]
  wire  _GEN_616 = hit_0 ? _GEN_104 : _GEN_488; // @[Cache_Soc.scala 96:19]
  wire  _GEN_617 = hit_0 ? _GEN_105 : _GEN_489; // @[Cache_Soc.scala 96:19]
  wire  _GEN_618 = hit_0 ? _GEN_106 : _GEN_490; // @[Cache_Soc.scala 96:19]
  wire  _GEN_619 = hit_0 ? _GEN_107 : _GEN_491; // @[Cache_Soc.scala 96:19]
  wire  _GEN_620 = hit_0 ? _GEN_108 : _GEN_492; // @[Cache_Soc.scala 96:19]
  wire  _GEN_621 = hit_0 ? _GEN_109 : _GEN_493; // @[Cache_Soc.scala 96:19]
  wire  _GEN_622 = hit_0 ? _GEN_110 : _GEN_494; // @[Cache_Soc.scala 96:19]
  wire  _GEN_623 = hit_0 ? _GEN_111 : _GEN_495; // @[Cache_Soc.scala 96:19]
  wire  _GEN_624 = hit_0 ? _GEN_112 : _GEN_496; // @[Cache_Soc.scala 96:19]
  wire  _GEN_625 = hit_0 ? _GEN_113 : _GEN_497; // @[Cache_Soc.scala 96:19]
  wire  _GEN_626 = hit_0 ? _GEN_114 : _GEN_498; // @[Cache_Soc.scala 96:19]
  wire  _GEN_627 = hit_0 ? _GEN_115 : _GEN_499; // @[Cache_Soc.scala 96:19]
  wire  _GEN_628 = hit_0 ? _GEN_116 : _GEN_500; // @[Cache_Soc.scala 96:19]
  wire  _GEN_629 = hit_0 ? _GEN_117 : _GEN_501; // @[Cache_Soc.scala 96:19]
  wire  _GEN_630 = hit_0 ? _GEN_118 : _GEN_502; // @[Cache_Soc.scala 96:19]
  wire  _GEN_631 = hit_0 ? _GEN_119 : _GEN_503; // @[Cache_Soc.scala 96:19]
  wire  _GEN_632 = hit_0 ? _GEN_120 : _GEN_504; // @[Cache_Soc.scala 96:19]
  wire  _GEN_633 = hit_0 ? _GEN_121 : _GEN_505; // @[Cache_Soc.scala 96:19]
  wire  _GEN_634 = hit_0 ? _GEN_122 : _GEN_506; // @[Cache_Soc.scala 96:19]
  wire  _GEN_635 = hit_0 ? _GEN_123 : _GEN_507; // @[Cache_Soc.scala 96:19]
  wire  _GEN_636 = hit_0 ? _GEN_124 : _GEN_508; // @[Cache_Soc.scala 96:19]
  wire  _GEN_637 = hit_0 ? _GEN_125 : _GEN_509; // @[Cache_Soc.scala 96:19]
  wire  _GEN_638 = hit_0 ? _GEN_126 : _GEN_510; // @[Cache_Soc.scala 96:19]
  wire  _GEN_639 = hit_0 ? _GEN_127 : _GEN_511; // @[Cache_Soc.scala 96:19]
  wire  _GEN_640 = hit_0 ? plru2_0 : _GEN_512; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_641 = hit_0 ? plru2_1 : _GEN_513; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_642 = hit_0 ? plru2_2 : _GEN_514; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_643 = hit_0 ? plru2_3 : _GEN_515; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_644 = hit_0 ? plru2_4 : _GEN_516; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_645 = hit_0 ? plru2_5 : _GEN_517; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_646 = hit_0 ? plru2_6 : _GEN_518; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_647 = hit_0 ? plru2_7 : _GEN_519; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_648 = hit_0 ? plru2_8 : _GEN_520; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_649 = hit_0 ? plru2_9 : _GEN_521; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_650 = hit_0 ? plru2_10 : _GEN_522; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_651 = hit_0 ? plru2_11 : _GEN_523; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_652 = hit_0 ? plru2_12 : _GEN_524; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_653 = hit_0 ? plru2_13 : _GEN_525; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_654 = hit_0 ? plru2_14 : _GEN_526; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_655 = hit_0 ? plru2_15 : _GEN_527; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_656 = hit_0 ? plru2_16 : _GEN_528; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_657 = hit_0 ? plru2_17 : _GEN_529; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_658 = hit_0 ? plru2_18 : _GEN_530; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_659 = hit_0 ? plru2_19 : _GEN_531; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_660 = hit_0 ? plru2_20 : _GEN_532; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_661 = hit_0 ? plru2_21 : _GEN_533; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_662 = hit_0 ? plru2_22 : _GEN_534; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_663 = hit_0 ? plru2_23 : _GEN_535; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_664 = hit_0 ? plru2_24 : _GEN_536; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_665 = hit_0 ? plru2_25 : _GEN_537; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_666 = hit_0 ? plru2_26 : _GEN_538; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_667 = hit_0 ? plru2_27 : _GEN_539; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_668 = hit_0 ? plru2_28 : _GEN_540; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_669 = hit_0 ? plru2_29 : _GEN_541; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_670 = hit_0 ? plru2_30 : _GEN_542; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_671 = hit_0 ? plru2_31 : _GEN_543; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_672 = hit_0 ? plru2_32 : _GEN_544; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_673 = hit_0 ? plru2_33 : _GEN_545; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_674 = hit_0 ? plru2_34 : _GEN_546; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_675 = hit_0 ? plru2_35 : _GEN_547; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_676 = hit_0 ? plru2_36 : _GEN_548; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_677 = hit_0 ? plru2_37 : _GEN_549; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_678 = hit_0 ? plru2_38 : _GEN_550; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_679 = hit_0 ? plru2_39 : _GEN_551; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_680 = hit_0 ? plru2_40 : _GEN_552; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_681 = hit_0 ? plru2_41 : _GEN_553; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_682 = hit_0 ? plru2_42 : _GEN_554; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_683 = hit_0 ? plru2_43 : _GEN_555; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_684 = hit_0 ? plru2_44 : _GEN_556; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_685 = hit_0 ? plru2_45 : _GEN_557; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_686 = hit_0 ? plru2_46 : _GEN_558; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_687 = hit_0 ? plru2_47 : _GEN_559; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_688 = hit_0 ? plru2_48 : _GEN_560; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_689 = hit_0 ? plru2_49 : _GEN_561; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_690 = hit_0 ? plru2_50 : _GEN_562; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_691 = hit_0 ? plru2_51 : _GEN_563; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_692 = hit_0 ? plru2_52 : _GEN_564; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_693 = hit_0 ? plru2_53 : _GEN_565; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_694 = hit_0 ? plru2_54 : _GEN_566; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_695 = hit_0 ? plru2_55 : _GEN_567; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_696 = hit_0 ? plru2_56 : _GEN_568; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_697 = hit_0 ? plru2_57 : _GEN_569; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_698 = hit_0 ? plru2_58 : _GEN_570; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_699 = hit_0 ? plru2_59 : _GEN_571; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_700 = hit_0 ? plru2_60 : _GEN_572; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_701 = hit_0 ? plru2_61 : _GEN_573; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_702 = hit_0 ? plru2_62 : _GEN_574; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_703 = hit_0 ? plru2_63 : _GEN_575; // @[Cache_Soc.scala 96:19 Cache_Soc.scala 91:22]
  wire  _GEN_704 = state == 3'h1 & cache_hit ? _GEN_0 : plru0_0; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_705 = state == 3'h1 & cache_hit ? _GEN_1 : plru0_1; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_706 = state == 3'h1 & cache_hit ? _GEN_2 : plru0_2; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_707 = state == 3'h1 & cache_hit ? _GEN_3 : plru0_3; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_708 = state == 3'h1 & cache_hit ? _GEN_4 : plru0_4; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_709 = state == 3'h1 & cache_hit ? _GEN_5 : plru0_5; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_710 = state == 3'h1 & cache_hit ? _GEN_6 : plru0_6; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_711 = state == 3'h1 & cache_hit ? _GEN_7 : plru0_7; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_712 = state == 3'h1 & cache_hit ? _GEN_8 : plru0_8; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_713 = state == 3'h1 & cache_hit ? _GEN_9 : plru0_9; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_714 = state == 3'h1 & cache_hit ? _GEN_10 : plru0_10; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_715 = state == 3'h1 & cache_hit ? _GEN_11 : plru0_11; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_716 = state == 3'h1 & cache_hit ? _GEN_12 : plru0_12; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_717 = state == 3'h1 & cache_hit ? _GEN_13 : plru0_13; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_718 = state == 3'h1 & cache_hit ? _GEN_14 : plru0_14; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_719 = state == 3'h1 & cache_hit ? _GEN_15 : plru0_15; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_720 = state == 3'h1 & cache_hit ? _GEN_16 : plru0_16; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_721 = state == 3'h1 & cache_hit ? _GEN_17 : plru0_17; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_722 = state == 3'h1 & cache_hit ? _GEN_18 : plru0_18; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_723 = state == 3'h1 & cache_hit ? _GEN_19 : plru0_19; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_724 = state == 3'h1 & cache_hit ? _GEN_20 : plru0_20; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_725 = state == 3'h1 & cache_hit ? _GEN_21 : plru0_21; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_726 = state == 3'h1 & cache_hit ? _GEN_22 : plru0_22; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_727 = state == 3'h1 & cache_hit ? _GEN_23 : plru0_23; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_728 = state == 3'h1 & cache_hit ? _GEN_24 : plru0_24; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_729 = state == 3'h1 & cache_hit ? _GEN_25 : plru0_25; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_730 = state == 3'h1 & cache_hit ? _GEN_26 : plru0_26; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_731 = state == 3'h1 & cache_hit ? _GEN_27 : plru0_27; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_732 = state == 3'h1 & cache_hit ? _GEN_28 : plru0_28; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_733 = state == 3'h1 & cache_hit ? _GEN_29 : plru0_29; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_734 = state == 3'h1 & cache_hit ? _GEN_30 : plru0_30; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_735 = state == 3'h1 & cache_hit ? _GEN_31 : plru0_31; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_736 = state == 3'h1 & cache_hit ? _GEN_32 : plru0_32; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_737 = state == 3'h1 & cache_hit ? _GEN_33 : plru0_33; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_738 = state == 3'h1 & cache_hit ? _GEN_34 : plru0_34; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_739 = state == 3'h1 & cache_hit ? _GEN_35 : plru0_35; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_740 = state == 3'h1 & cache_hit ? _GEN_36 : plru0_36; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_741 = state == 3'h1 & cache_hit ? _GEN_37 : plru0_37; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_742 = state == 3'h1 & cache_hit ? _GEN_38 : plru0_38; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_743 = state == 3'h1 & cache_hit ? _GEN_39 : plru0_39; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_744 = state == 3'h1 & cache_hit ? _GEN_40 : plru0_40; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_745 = state == 3'h1 & cache_hit ? _GEN_41 : plru0_41; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_746 = state == 3'h1 & cache_hit ? _GEN_42 : plru0_42; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_747 = state == 3'h1 & cache_hit ? _GEN_43 : plru0_43; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_748 = state == 3'h1 & cache_hit ? _GEN_44 : plru0_44; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_749 = state == 3'h1 & cache_hit ? _GEN_45 : plru0_45; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_750 = state == 3'h1 & cache_hit ? _GEN_46 : plru0_46; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_751 = state == 3'h1 & cache_hit ? _GEN_47 : plru0_47; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_752 = state == 3'h1 & cache_hit ? _GEN_48 : plru0_48; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_753 = state == 3'h1 & cache_hit ? _GEN_49 : plru0_49; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_754 = state == 3'h1 & cache_hit ? _GEN_50 : plru0_50; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_755 = state == 3'h1 & cache_hit ? _GEN_51 : plru0_51; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_756 = state == 3'h1 & cache_hit ? _GEN_52 : plru0_52; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_757 = state == 3'h1 & cache_hit ? _GEN_53 : plru0_53; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_758 = state == 3'h1 & cache_hit ? _GEN_54 : plru0_54; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_759 = state == 3'h1 & cache_hit ? _GEN_55 : plru0_55; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_760 = state == 3'h1 & cache_hit ? _GEN_56 : plru0_56; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_761 = state == 3'h1 & cache_hit ? _GEN_57 : plru0_57; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_762 = state == 3'h1 & cache_hit ? _GEN_58 : plru0_58; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_763 = state == 3'h1 & cache_hit ? _GEN_59 : plru0_59; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_764 = state == 3'h1 & cache_hit ? _GEN_60 : plru0_60; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_765 = state == 3'h1 & cache_hit ? _GEN_61 : plru0_61; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_766 = state == 3'h1 & cache_hit ? _GEN_62 : plru0_62; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_767 = state == 3'h1 & cache_hit ? _GEN_63 : plru0_63; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 89:22]
  wire  _GEN_768 = state == 3'h1 & cache_hit ? _GEN_576 : plru1_0; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_769 = state == 3'h1 & cache_hit ? _GEN_577 : plru1_1; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_770 = state == 3'h1 & cache_hit ? _GEN_578 : plru1_2; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_771 = state == 3'h1 & cache_hit ? _GEN_579 : plru1_3; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_772 = state == 3'h1 & cache_hit ? _GEN_580 : plru1_4; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_773 = state == 3'h1 & cache_hit ? _GEN_581 : plru1_5; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_774 = state == 3'h1 & cache_hit ? _GEN_582 : plru1_6; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_775 = state == 3'h1 & cache_hit ? _GEN_583 : plru1_7; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_776 = state == 3'h1 & cache_hit ? _GEN_584 : plru1_8; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_777 = state == 3'h1 & cache_hit ? _GEN_585 : plru1_9; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_778 = state == 3'h1 & cache_hit ? _GEN_586 : plru1_10; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_779 = state == 3'h1 & cache_hit ? _GEN_587 : plru1_11; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_780 = state == 3'h1 & cache_hit ? _GEN_588 : plru1_12; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_781 = state == 3'h1 & cache_hit ? _GEN_589 : plru1_13; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_782 = state == 3'h1 & cache_hit ? _GEN_590 : plru1_14; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_783 = state == 3'h1 & cache_hit ? _GEN_591 : plru1_15; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_784 = state == 3'h1 & cache_hit ? _GEN_592 : plru1_16; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_785 = state == 3'h1 & cache_hit ? _GEN_593 : plru1_17; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_786 = state == 3'h1 & cache_hit ? _GEN_594 : plru1_18; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_787 = state == 3'h1 & cache_hit ? _GEN_595 : plru1_19; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_788 = state == 3'h1 & cache_hit ? _GEN_596 : plru1_20; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_789 = state == 3'h1 & cache_hit ? _GEN_597 : plru1_21; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_790 = state == 3'h1 & cache_hit ? _GEN_598 : plru1_22; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_791 = state == 3'h1 & cache_hit ? _GEN_599 : plru1_23; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_792 = state == 3'h1 & cache_hit ? _GEN_600 : plru1_24; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_793 = state == 3'h1 & cache_hit ? _GEN_601 : plru1_25; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_794 = state == 3'h1 & cache_hit ? _GEN_602 : plru1_26; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_795 = state == 3'h1 & cache_hit ? _GEN_603 : plru1_27; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_796 = state == 3'h1 & cache_hit ? _GEN_604 : plru1_28; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_797 = state == 3'h1 & cache_hit ? _GEN_605 : plru1_29; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_798 = state == 3'h1 & cache_hit ? _GEN_606 : plru1_30; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_799 = state == 3'h1 & cache_hit ? _GEN_607 : plru1_31; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_800 = state == 3'h1 & cache_hit ? _GEN_608 : plru1_32; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_801 = state == 3'h1 & cache_hit ? _GEN_609 : plru1_33; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_802 = state == 3'h1 & cache_hit ? _GEN_610 : plru1_34; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_803 = state == 3'h1 & cache_hit ? _GEN_611 : plru1_35; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_804 = state == 3'h1 & cache_hit ? _GEN_612 : plru1_36; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_805 = state == 3'h1 & cache_hit ? _GEN_613 : plru1_37; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_806 = state == 3'h1 & cache_hit ? _GEN_614 : plru1_38; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_807 = state == 3'h1 & cache_hit ? _GEN_615 : plru1_39; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_808 = state == 3'h1 & cache_hit ? _GEN_616 : plru1_40; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_809 = state == 3'h1 & cache_hit ? _GEN_617 : plru1_41; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_810 = state == 3'h1 & cache_hit ? _GEN_618 : plru1_42; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_811 = state == 3'h1 & cache_hit ? _GEN_619 : plru1_43; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_812 = state == 3'h1 & cache_hit ? _GEN_620 : plru1_44; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_813 = state == 3'h1 & cache_hit ? _GEN_621 : plru1_45; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_814 = state == 3'h1 & cache_hit ? _GEN_622 : plru1_46; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_815 = state == 3'h1 & cache_hit ? _GEN_623 : plru1_47; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_816 = state == 3'h1 & cache_hit ? _GEN_624 : plru1_48; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_817 = state == 3'h1 & cache_hit ? _GEN_625 : plru1_49; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_818 = state == 3'h1 & cache_hit ? _GEN_626 : plru1_50; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_819 = state == 3'h1 & cache_hit ? _GEN_627 : plru1_51; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_820 = state == 3'h1 & cache_hit ? _GEN_628 : plru1_52; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_821 = state == 3'h1 & cache_hit ? _GEN_629 : plru1_53; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_822 = state == 3'h1 & cache_hit ? _GEN_630 : plru1_54; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_823 = state == 3'h1 & cache_hit ? _GEN_631 : plru1_55; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_824 = state == 3'h1 & cache_hit ? _GEN_632 : plru1_56; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_825 = state == 3'h1 & cache_hit ? _GEN_633 : plru1_57; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_826 = state == 3'h1 & cache_hit ? _GEN_634 : plru1_58; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_827 = state == 3'h1 & cache_hit ? _GEN_635 : plru1_59; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_828 = state == 3'h1 & cache_hit ? _GEN_636 : plru1_60; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_829 = state == 3'h1 & cache_hit ? _GEN_637 : plru1_61; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_830 = state == 3'h1 & cache_hit ? _GEN_638 : plru1_62; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_831 = state == 3'h1 & cache_hit ? _GEN_639 : plru1_63; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 90:22]
  wire  _GEN_832 = state == 3'h1 & cache_hit ? _GEN_640 : plru2_0; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_833 = state == 3'h1 & cache_hit ? _GEN_641 : plru2_1; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_834 = state == 3'h1 & cache_hit ? _GEN_642 : plru2_2; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_835 = state == 3'h1 & cache_hit ? _GEN_643 : plru2_3; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_836 = state == 3'h1 & cache_hit ? _GEN_644 : plru2_4; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_837 = state == 3'h1 & cache_hit ? _GEN_645 : plru2_5; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_838 = state == 3'h1 & cache_hit ? _GEN_646 : plru2_6; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_839 = state == 3'h1 & cache_hit ? _GEN_647 : plru2_7; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_840 = state == 3'h1 & cache_hit ? _GEN_648 : plru2_8; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_841 = state == 3'h1 & cache_hit ? _GEN_649 : plru2_9; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_842 = state == 3'h1 & cache_hit ? _GEN_650 : plru2_10; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_843 = state == 3'h1 & cache_hit ? _GEN_651 : plru2_11; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_844 = state == 3'h1 & cache_hit ? _GEN_652 : plru2_12; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_845 = state == 3'h1 & cache_hit ? _GEN_653 : plru2_13; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_846 = state == 3'h1 & cache_hit ? _GEN_654 : plru2_14; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_847 = state == 3'h1 & cache_hit ? _GEN_655 : plru2_15; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_848 = state == 3'h1 & cache_hit ? _GEN_656 : plru2_16; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_849 = state == 3'h1 & cache_hit ? _GEN_657 : plru2_17; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_850 = state == 3'h1 & cache_hit ? _GEN_658 : plru2_18; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_851 = state == 3'h1 & cache_hit ? _GEN_659 : plru2_19; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_852 = state == 3'h1 & cache_hit ? _GEN_660 : plru2_20; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_853 = state == 3'h1 & cache_hit ? _GEN_661 : plru2_21; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_854 = state == 3'h1 & cache_hit ? _GEN_662 : plru2_22; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_855 = state == 3'h1 & cache_hit ? _GEN_663 : plru2_23; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_856 = state == 3'h1 & cache_hit ? _GEN_664 : plru2_24; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_857 = state == 3'h1 & cache_hit ? _GEN_665 : plru2_25; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_858 = state == 3'h1 & cache_hit ? _GEN_666 : plru2_26; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_859 = state == 3'h1 & cache_hit ? _GEN_667 : plru2_27; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_860 = state == 3'h1 & cache_hit ? _GEN_668 : plru2_28; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_861 = state == 3'h1 & cache_hit ? _GEN_669 : plru2_29; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_862 = state == 3'h1 & cache_hit ? _GEN_670 : plru2_30; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_863 = state == 3'h1 & cache_hit ? _GEN_671 : plru2_31; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_864 = state == 3'h1 & cache_hit ? _GEN_672 : plru2_32; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_865 = state == 3'h1 & cache_hit ? _GEN_673 : plru2_33; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_866 = state == 3'h1 & cache_hit ? _GEN_674 : plru2_34; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_867 = state == 3'h1 & cache_hit ? _GEN_675 : plru2_35; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_868 = state == 3'h1 & cache_hit ? _GEN_676 : plru2_36; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_869 = state == 3'h1 & cache_hit ? _GEN_677 : plru2_37; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_870 = state == 3'h1 & cache_hit ? _GEN_678 : plru2_38; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_871 = state == 3'h1 & cache_hit ? _GEN_679 : plru2_39; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_872 = state == 3'h1 & cache_hit ? _GEN_680 : plru2_40; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_873 = state == 3'h1 & cache_hit ? _GEN_681 : plru2_41; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_874 = state == 3'h1 & cache_hit ? _GEN_682 : plru2_42; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_875 = state == 3'h1 & cache_hit ? _GEN_683 : plru2_43; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_876 = state == 3'h1 & cache_hit ? _GEN_684 : plru2_44; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_877 = state == 3'h1 & cache_hit ? _GEN_685 : plru2_45; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_878 = state == 3'h1 & cache_hit ? _GEN_686 : plru2_46; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_879 = state == 3'h1 & cache_hit ? _GEN_687 : plru2_47; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_880 = state == 3'h1 & cache_hit ? _GEN_688 : plru2_48; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_881 = state == 3'h1 & cache_hit ? _GEN_689 : plru2_49; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_882 = state == 3'h1 & cache_hit ? _GEN_690 : plru2_50; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_883 = state == 3'h1 & cache_hit ? _GEN_691 : plru2_51; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_884 = state == 3'h1 & cache_hit ? _GEN_692 : plru2_52; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_885 = state == 3'h1 & cache_hit ? _GEN_693 : plru2_53; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_886 = state == 3'h1 & cache_hit ? _GEN_694 : plru2_54; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_887 = state == 3'h1 & cache_hit ? _GEN_695 : plru2_55; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_888 = state == 3'h1 & cache_hit ? _GEN_696 : plru2_56; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_889 = state == 3'h1 & cache_hit ? _GEN_697 : plru2_57; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_890 = state == 3'h1 & cache_hit ? _GEN_698 : plru2_58; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_891 = state == 3'h1 & cache_hit ? _GEN_699 : plru2_59; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_892 = state == 3'h1 & cache_hit ? _GEN_700 : plru2_60; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_893 = state == 3'h1 & cache_hit ? _GEN_701 : plru2_61; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_894 = state == 3'h1 & cache_hit ? _GEN_702 : plru2_62; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _GEN_895 = state == 3'h1 & cache_hit ? _GEN_703 : plru2_63; // @[Cache_Soc.scala 94:42 Cache_Soc.scala 91:22]
  wire  _T_2 = state == 3'h4; // @[Cache_Soc.scala 106:16]
  wire  _T_3 = state == 3'h4 & io_out_ret_valid; // @[Cache_Soc.scala 106:28]
  wire  _GEN_1793 = 6'h1 == rb_index ? plru0_1 : plru0_0; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1794 = 6'h2 == rb_index ? plru0_2 : _GEN_1793; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1795 = 6'h3 == rb_index ? plru0_3 : _GEN_1794; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1796 = 6'h4 == rb_index ? plru0_4 : _GEN_1795; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1797 = 6'h5 == rb_index ? plru0_5 : _GEN_1796; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1798 = 6'h6 == rb_index ? plru0_6 : _GEN_1797; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1799 = 6'h7 == rb_index ? plru0_7 : _GEN_1798; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1800 = 6'h8 == rb_index ? plru0_8 : _GEN_1799; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1801 = 6'h9 == rb_index ? plru0_9 : _GEN_1800; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1802 = 6'ha == rb_index ? plru0_10 : _GEN_1801; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1803 = 6'hb == rb_index ? plru0_11 : _GEN_1802; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1804 = 6'hc == rb_index ? plru0_12 : _GEN_1803; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1805 = 6'hd == rb_index ? plru0_13 : _GEN_1804; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1806 = 6'he == rb_index ? plru0_14 : _GEN_1805; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1807 = 6'hf == rb_index ? plru0_15 : _GEN_1806; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1808 = 6'h10 == rb_index ? plru0_16 : _GEN_1807; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1809 = 6'h11 == rb_index ? plru0_17 : _GEN_1808; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1810 = 6'h12 == rb_index ? plru0_18 : _GEN_1809; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1811 = 6'h13 == rb_index ? plru0_19 : _GEN_1810; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1812 = 6'h14 == rb_index ? plru0_20 : _GEN_1811; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1813 = 6'h15 == rb_index ? plru0_21 : _GEN_1812; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1814 = 6'h16 == rb_index ? plru0_22 : _GEN_1813; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1815 = 6'h17 == rb_index ? plru0_23 : _GEN_1814; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1816 = 6'h18 == rb_index ? plru0_24 : _GEN_1815; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1817 = 6'h19 == rb_index ? plru0_25 : _GEN_1816; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1818 = 6'h1a == rb_index ? plru0_26 : _GEN_1817; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1819 = 6'h1b == rb_index ? plru0_27 : _GEN_1818; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1820 = 6'h1c == rb_index ? plru0_28 : _GEN_1819; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1821 = 6'h1d == rb_index ? plru0_29 : _GEN_1820; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1822 = 6'h1e == rb_index ? plru0_30 : _GEN_1821; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1823 = 6'h1f == rb_index ? plru0_31 : _GEN_1822; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1824 = 6'h20 == rb_index ? plru0_32 : _GEN_1823; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1825 = 6'h21 == rb_index ? plru0_33 : _GEN_1824; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1826 = 6'h22 == rb_index ? plru0_34 : _GEN_1825; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1827 = 6'h23 == rb_index ? plru0_35 : _GEN_1826; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1828 = 6'h24 == rb_index ? plru0_36 : _GEN_1827; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1829 = 6'h25 == rb_index ? plru0_37 : _GEN_1828; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1830 = 6'h26 == rb_index ? plru0_38 : _GEN_1829; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1831 = 6'h27 == rb_index ? plru0_39 : _GEN_1830; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1832 = 6'h28 == rb_index ? plru0_40 : _GEN_1831; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1833 = 6'h29 == rb_index ? plru0_41 : _GEN_1832; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1834 = 6'h2a == rb_index ? plru0_42 : _GEN_1833; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1835 = 6'h2b == rb_index ? plru0_43 : _GEN_1834; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1836 = 6'h2c == rb_index ? plru0_44 : _GEN_1835; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1837 = 6'h2d == rb_index ? plru0_45 : _GEN_1836; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1838 = 6'h2e == rb_index ? plru0_46 : _GEN_1837; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1839 = 6'h2f == rb_index ? plru0_47 : _GEN_1838; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1840 = 6'h30 == rb_index ? plru0_48 : _GEN_1839; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1841 = 6'h31 == rb_index ? plru0_49 : _GEN_1840; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1842 = 6'h32 == rb_index ? plru0_50 : _GEN_1841; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1843 = 6'h33 == rb_index ? plru0_51 : _GEN_1842; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1844 = 6'h34 == rb_index ? plru0_52 : _GEN_1843; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1845 = 6'h35 == rb_index ? plru0_53 : _GEN_1844; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1846 = 6'h36 == rb_index ? plru0_54 : _GEN_1845; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1847 = 6'h37 == rb_index ? plru0_55 : _GEN_1846; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1848 = 6'h38 == rb_index ? plru0_56 : _GEN_1847; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1849 = 6'h39 == rb_index ? plru0_57 : _GEN_1848; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1850 = 6'h3a == rb_index ? plru0_58 : _GEN_1849; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1851 = 6'h3b == rb_index ? plru0_59 : _GEN_1850; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1852 = 6'h3c == rb_index ? plru0_60 : _GEN_1851; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1853 = 6'h3d == rb_index ? plru0_61 : _GEN_1852; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1854 = 6'h3e == rb_index ? plru0_62 : _GEN_1853; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1855 = 6'h3f == rb_index ? plru0_63 : _GEN_1854; // @[Cache_Soc.scala 119:59 Cache_Soc.scala 119:59]
  wire  _GEN_1857 = 6'h1 == rb_index ? plru1_1 : plru1_0; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1858 = 6'h2 == rb_index ? plru1_2 : _GEN_1857; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1859 = 6'h3 == rb_index ? plru1_3 : _GEN_1858; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1860 = 6'h4 == rb_index ? plru1_4 : _GEN_1859; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1861 = 6'h5 == rb_index ? plru1_5 : _GEN_1860; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1862 = 6'h6 == rb_index ? plru1_6 : _GEN_1861; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1863 = 6'h7 == rb_index ? plru1_7 : _GEN_1862; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1864 = 6'h8 == rb_index ? plru1_8 : _GEN_1863; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1865 = 6'h9 == rb_index ? plru1_9 : _GEN_1864; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1866 = 6'ha == rb_index ? plru1_10 : _GEN_1865; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1867 = 6'hb == rb_index ? plru1_11 : _GEN_1866; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1868 = 6'hc == rb_index ? plru1_12 : _GEN_1867; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1869 = 6'hd == rb_index ? plru1_13 : _GEN_1868; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1870 = 6'he == rb_index ? plru1_14 : _GEN_1869; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1871 = 6'hf == rb_index ? plru1_15 : _GEN_1870; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1872 = 6'h10 == rb_index ? plru1_16 : _GEN_1871; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1873 = 6'h11 == rb_index ? plru1_17 : _GEN_1872; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1874 = 6'h12 == rb_index ? plru1_18 : _GEN_1873; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1875 = 6'h13 == rb_index ? plru1_19 : _GEN_1874; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1876 = 6'h14 == rb_index ? plru1_20 : _GEN_1875; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1877 = 6'h15 == rb_index ? plru1_21 : _GEN_1876; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1878 = 6'h16 == rb_index ? plru1_22 : _GEN_1877; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1879 = 6'h17 == rb_index ? plru1_23 : _GEN_1878; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1880 = 6'h18 == rb_index ? plru1_24 : _GEN_1879; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1881 = 6'h19 == rb_index ? plru1_25 : _GEN_1880; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1882 = 6'h1a == rb_index ? plru1_26 : _GEN_1881; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1883 = 6'h1b == rb_index ? plru1_27 : _GEN_1882; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1884 = 6'h1c == rb_index ? plru1_28 : _GEN_1883; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1885 = 6'h1d == rb_index ? plru1_29 : _GEN_1884; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1886 = 6'h1e == rb_index ? plru1_30 : _GEN_1885; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1887 = 6'h1f == rb_index ? plru1_31 : _GEN_1886; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1888 = 6'h20 == rb_index ? plru1_32 : _GEN_1887; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1889 = 6'h21 == rb_index ? plru1_33 : _GEN_1888; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1890 = 6'h22 == rb_index ? plru1_34 : _GEN_1889; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1891 = 6'h23 == rb_index ? plru1_35 : _GEN_1890; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1892 = 6'h24 == rb_index ? plru1_36 : _GEN_1891; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1893 = 6'h25 == rb_index ? plru1_37 : _GEN_1892; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1894 = 6'h26 == rb_index ? plru1_38 : _GEN_1893; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1895 = 6'h27 == rb_index ? plru1_39 : _GEN_1894; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1896 = 6'h28 == rb_index ? plru1_40 : _GEN_1895; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1897 = 6'h29 == rb_index ? plru1_41 : _GEN_1896; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1898 = 6'h2a == rb_index ? plru1_42 : _GEN_1897; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1899 = 6'h2b == rb_index ? plru1_43 : _GEN_1898; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1900 = 6'h2c == rb_index ? plru1_44 : _GEN_1899; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1901 = 6'h2d == rb_index ? plru1_45 : _GEN_1900; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1902 = 6'h2e == rb_index ? plru1_46 : _GEN_1901; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1903 = 6'h2f == rb_index ? plru1_47 : _GEN_1902; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1904 = 6'h30 == rb_index ? plru1_48 : _GEN_1903; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1905 = 6'h31 == rb_index ? plru1_49 : _GEN_1904; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1906 = 6'h32 == rb_index ? plru1_50 : _GEN_1905; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1907 = 6'h33 == rb_index ? plru1_51 : _GEN_1906; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1908 = 6'h34 == rb_index ? plru1_52 : _GEN_1907; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1909 = 6'h35 == rb_index ? plru1_53 : _GEN_1908; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1910 = 6'h36 == rb_index ? plru1_54 : _GEN_1909; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1911 = 6'h37 == rb_index ? plru1_55 : _GEN_1910; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1912 = 6'h38 == rb_index ? plru1_56 : _GEN_1911; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1913 = 6'h39 == rb_index ? plru1_57 : _GEN_1912; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1914 = 6'h3a == rb_index ? plru1_58 : _GEN_1913; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1915 = 6'h3b == rb_index ? plru1_59 : _GEN_1914; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1916 = 6'h3c == rb_index ? plru1_60 : _GEN_1915; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1917 = 6'h3d == rb_index ? plru1_61 : _GEN_1916; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1918 = 6'h3e == rb_index ? plru1_62 : _GEN_1917; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1919 = 6'h3f == rb_index ? plru1_63 : _GEN_1918; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1921 = 6'h1 == rb_index ? plru2_1 : plru2_0; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1922 = 6'h2 == rb_index ? plru2_2 : _GEN_1921; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1923 = 6'h3 == rb_index ? plru2_3 : _GEN_1922; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1924 = 6'h4 == rb_index ? plru2_4 : _GEN_1923; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1925 = 6'h5 == rb_index ? plru2_5 : _GEN_1924; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1926 = 6'h6 == rb_index ? plru2_6 : _GEN_1925; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1927 = 6'h7 == rb_index ? plru2_7 : _GEN_1926; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1928 = 6'h8 == rb_index ? plru2_8 : _GEN_1927; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1929 = 6'h9 == rb_index ? plru2_9 : _GEN_1928; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1930 = 6'ha == rb_index ? plru2_10 : _GEN_1929; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1931 = 6'hb == rb_index ? plru2_11 : _GEN_1930; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1932 = 6'hc == rb_index ? plru2_12 : _GEN_1931; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1933 = 6'hd == rb_index ? plru2_13 : _GEN_1932; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1934 = 6'he == rb_index ? plru2_14 : _GEN_1933; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1935 = 6'hf == rb_index ? plru2_15 : _GEN_1934; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1936 = 6'h10 == rb_index ? plru2_16 : _GEN_1935; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1937 = 6'h11 == rb_index ? plru2_17 : _GEN_1936; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1938 = 6'h12 == rb_index ? plru2_18 : _GEN_1937; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1939 = 6'h13 == rb_index ? plru2_19 : _GEN_1938; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1940 = 6'h14 == rb_index ? plru2_20 : _GEN_1939; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1941 = 6'h15 == rb_index ? plru2_21 : _GEN_1940; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1942 = 6'h16 == rb_index ? plru2_22 : _GEN_1941; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1943 = 6'h17 == rb_index ? plru2_23 : _GEN_1942; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1944 = 6'h18 == rb_index ? plru2_24 : _GEN_1943; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1945 = 6'h19 == rb_index ? plru2_25 : _GEN_1944; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1946 = 6'h1a == rb_index ? plru2_26 : _GEN_1945; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1947 = 6'h1b == rb_index ? plru2_27 : _GEN_1946; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1948 = 6'h1c == rb_index ? plru2_28 : _GEN_1947; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1949 = 6'h1d == rb_index ? plru2_29 : _GEN_1948; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1950 = 6'h1e == rb_index ? plru2_30 : _GEN_1949; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1951 = 6'h1f == rb_index ? plru2_31 : _GEN_1950; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1952 = 6'h20 == rb_index ? plru2_32 : _GEN_1951; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1953 = 6'h21 == rb_index ? plru2_33 : _GEN_1952; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1954 = 6'h22 == rb_index ? plru2_34 : _GEN_1953; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1955 = 6'h23 == rb_index ? plru2_35 : _GEN_1954; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1956 = 6'h24 == rb_index ? plru2_36 : _GEN_1955; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1957 = 6'h25 == rb_index ? plru2_37 : _GEN_1956; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1958 = 6'h26 == rb_index ? plru2_38 : _GEN_1957; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1959 = 6'h27 == rb_index ? plru2_39 : _GEN_1958; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1960 = 6'h28 == rb_index ? plru2_40 : _GEN_1959; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1961 = 6'h29 == rb_index ? plru2_41 : _GEN_1960; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1962 = 6'h2a == rb_index ? plru2_42 : _GEN_1961; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1963 = 6'h2b == rb_index ? plru2_43 : _GEN_1962; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1964 = 6'h2c == rb_index ? plru2_44 : _GEN_1963; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1965 = 6'h2d == rb_index ? plru2_45 : _GEN_1964; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1966 = 6'h2e == rb_index ? plru2_46 : _GEN_1965; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1967 = 6'h2f == rb_index ? plru2_47 : _GEN_1966; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1968 = 6'h30 == rb_index ? plru2_48 : _GEN_1967; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1969 = 6'h31 == rb_index ? plru2_49 : _GEN_1968; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1970 = 6'h32 == rb_index ? plru2_50 : _GEN_1969; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1971 = 6'h33 == rb_index ? plru2_51 : _GEN_1970; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1972 = 6'h34 == rb_index ? plru2_52 : _GEN_1971; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1973 = 6'h35 == rb_index ? plru2_53 : _GEN_1972; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1974 = 6'h36 == rb_index ? plru2_54 : _GEN_1973; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1975 = 6'h37 == rb_index ? plru2_55 : _GEN_1974; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1976 = 6'h38 == rb_index ? plru2_56 : _GEN_1975; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1977 = 6'h39 == rb_index ? plru2_57 : _GEN_1976; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1978 = 6'h3a == rb_index ? plru2_58 : _GEN_1977; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1979 = 6'h3b == rb_index ? plru2_59 : _GEN_1978; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1980 = 6'h3c == rb_index ? plru2_60 : _GEN_1979; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1981 = 6'h3d == rb_index ? plru2_61 : _GEN_1980; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1982 = 6'h3e == rb_index ? plru2_62 : _GEN_1981; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  _GEN_1983 = 6'h3f == rb_index ? plru2_63 : _GEN_1982; // @[Cache_Soc.scala 119:42 Cache_Soc.scala 119:42]
  wire  replace_way_lo = ~_GEN_1855 ? _GEN_1919 : _GEN_1983; // @[Cache_Soc.scala 119:42]
  wire [1:0] replace_way = {_GEN_1855,replace_way_lo}; // @[Cat.scala 30:58]
  wire  _plru0_T_1 = replace_way == 2'h0; // @[Cache_Soc.scala 107:36]
  wire  _plru0_T_2 = replace_way == 2'h1; // @[Cache_Soc.scala 107:59]
  wire  _GEN_960 = _GEN_2439 | _GEN_768; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_961 = _GEN_2440 | _GEN_769; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_962 = _GEN_2441 | _GEN_770; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_963 = _GEN_2442 | _GEN_771; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_964 = _GEN_2443 | _GEN_772; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_965 = _GEN_2444 | _GEN_773; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_966 = _GEN_2445 | _GEN_774; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_967 = _GEN_2446 | _GEN_775; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_968 = _GEN_2447 | _GEN_776; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_969 = _GEN_2448 | _GEN_777; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_970 = _GEN_2449 | _GEN_778; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_971 = _GEN_2450 | _GEN_779; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_972 = _GEN_2451 | _GEN_780; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_973 = _GEN_2452 | _GEN_781; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_974 = _GEN_2453 | _GEN_782; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_975 = _GEN_2454 | _GEN_783; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_976 = _GEN_2455 | _GEN_784; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_977 = _GEN_2456 | _GEN_785; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_978 = _GEN_2457 | _GEN_786; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_979 = _GEN_2458 | _GEN_787; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_980 = _GEN_2459 | _GEN_788; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_981 = _GEN_2460 | _GEN_789; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_982 = _GEN_2461 | _GEN_790; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_983 = _GEN_2462 | _GEN_791; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_984 = _GEN_2463 | _GEN_792; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_985 = _GEN_2464 | _GEN_793; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_986 = _GEN_2465 | _GEN_794; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_987 = _GEN_2466 | _GEN_795; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_988 = _GEN_2467 | _GEN_796; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_989 = _GEN_2468 | _GEN_797; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_990 = _GEN_2469 | _GEN_798; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_991 = _GEN_2470 | _GEN_799; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_992 = _GEN_2471 | _GEN_800; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_993 = _GEN_2472 | _GEN_801; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_994 = _GEN_2473 | _GEN_802; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_995 = _GEN_2474 | _GEN_803; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_996 = _GEN_2475 | _GEN_804; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_997 = _GEN_2476 | _GEN_805; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_998 = _GEN_2477 | _GEN_806; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_999 = _GEN_2478 | _GEN_807; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1000 = _GEN_2479 | _GEN_808; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1001 = _GEN_2480 | _GEN_809; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1002 = _GEN_2481 | _GEN_810; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1003 = _GEN_2482 | _GEN_811; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1004 = _GEN_2483 | _GEN_812; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1005 = _GEN_2484 | _GEN_813; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1006 = _GEN_2485 | _GEN_814; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1007 = _GEN_2486 | _GEN_815; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1008 = _GEN_2487 | _GEN_816; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1009 = _GEN_2488 | _GEN_817; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1010 = _GEN_2489 | _GEN_818; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1011 = _GEN_2490 | _GEN_819; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1012 = _GEN_2491 | _GEN_820; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1013 = _GEN_2492 | _GEN_821; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1014 = _GEN_2493 | _GEN_822; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1015 = _GEN_2494 | _GEN_823; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1016 = _GEN_2495 | _GEN_824; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1017 = _GEN_2496 | _GEN_825; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1018 = _GEN_2497 | _GEN_826; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1019 = _GEN_2498 | _GEN_827; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1020 = _GEN_2499 | _GEN_828; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1021 = _GEN_2500 | _GEN_829; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1022 = _GEN_2501 | _GEN_830; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1023 = _GEN_2502 | _GEN_831; // @[Cache_Soc.scala 109:23 Cache_Soc.scala 109:23]
  wire  _GEN_1024 = 6'h0 == rb_index ? 1'h0 : _GEN_768; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1025 = 6'h1 == rb_index ? 1'h0 : _GEN_769; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1026 = 6'h2 == rb_index ? 1'h0 : _GEN_770; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1027 = 6'h3 == rb_index ? 1'h0 : _GEN_771; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1028 = 6'h4 == rb_index ? 1'h0 : _GEN_772; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1029 = 6'h5 == rb_index ? 1'h0 : _GEN_773; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1030 = 6'h6 == rb_index ? 1'h0 : _GEN_774; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1031 = 6'h7 == rb_index ? 1'h0 : _GEN_775; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1032 = 6'h8 == rb_index ? 1'h0 : _GEN_776; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1033 = 6'h9 == rb_index ? 1'h0 : _GEN_777; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1034 = 6'ha == rb_index ? 1'h0 : _GEN_778; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1035 = 6'hb == rb_index ? 1'h0 : _GEN_779; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1036 = 6'hc == rb_index ? 1'h0 : _GEN_780; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1037 = 6'hd == rb_index ? 1'h0 : _GEN_781; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1038 = 6'he == rb_index ? 1'h0 : _GEN_782; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1039 = 6'hf == rb_index ? 1'h0 : _GEN_783; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1040 = 6'h10 == rb_index ? 1'h0 : _GEN_784; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1041 = 6'h11 == rb_index ? 1'h0 : _GEN_785; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1042 = 6'h12 == rb_index ? 1'h0 : _GEN_786; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1043 = 6'h13 == rb_index ? 1'h0 : _GEN_787; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1044 = 6'h14 == rb_index ? 1'h0 : _GEN_788; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1045 = 6'h15 == rb_index ? 1'h0 : _GEN_789; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1046 = 6'h16 == rb_index ? 1'h0 : _GEN_790; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1047 = 6'h17 == rb_index ? 1'h0 : _GEN_791; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1048 = 6'h18 == rb_index ? 1'h0 : _GEN_792; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1049 = 6'h19 == rb_index ? 1'h0 : _GEN_793; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1050 = 6'h1a == rb_index ? 1'h0 : _GEN_794; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1051 = 6'h1b == rb_index ? 1'h0 : _GEN_795; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1052 = 6'h1c == rb_index ? 1'h0 : _GEN_796; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1053 = 6'h1d == rb_index ? 1'h0 : _GEN_797; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1054 = 6'h1e == rb_index ? 1'h0 : _GEN_798; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1055 = 6'h1f == rb_index ? 1'h0 : _GEN_799; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1056 = 6'h20 == rb_index ? 1'h0 : _GEN_800; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1057 = 6'h21 == rb_index ? 1'h0 : _GEN_801; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1058 = 6'h22 == rb_index ? 1'h0 : _GEN_802; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1059 = 6'h23 == rb_index ? 1'h0 : _GEN_803; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1060 = 6'h24 == rb_index ? 1'h0 : _GEN_804; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1061 = 6'h25 == rb_index ? 1'h0 : _GEN_805; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1062 = 6'h26 == rb_index ? 1'h0 : _GEN_806; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1063 = 6'h27 == rb_index ? 1'h0 : _GEN_807; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1064 = 6'h28 == rb_index ? 1'h0 : _GEN_808; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1065 = 6'h29 == rb_index ? 1'h0 : _GEN_809; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1066 = 6'h2a == rb_index ? 1'h0 : _GEN_810; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1067 = 6'h2b == rb_index ? 1'h0 : _GEN_811; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1068 = 6'h2c == rb_index ? 1'h0 : _GEN_812; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1069 = 6'h2d == rb_index ? 1'h0 : _GEN_813; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1070 = 6'h2e == rb_index ? 1'h0 : _GEN_814; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1071 = 6'h2f == rb_index ? 1'h0 : _GEN_815; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1072 = 6'h30 == rb_index ? 1'h0 : _GEN_816; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1073 = 6'h31 == rb_index ? 1'h0 : _GEN_817; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1074 = 6'h32 == rb_index ? 1'h0 : _GEN_818; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1075 = 6'h33 == rb_index ? 1'h0 : _GEN_819; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1076 = 6'h34 == rb_index ? 1'h0 : _GEN_820; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1077 = 6'h35 == rb_index ? 1'h0 : _GEN_821; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1078 = 6'h36 == rb_index ? 1'h0 : _GEN_822; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1079 = 6'h37 == rb_index ? 1'h0 : _GEN_823; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1080 = 6'h38 == rb_index ? 1'h0 : _GEN_824; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1081 = 6'h39 == rb_index ? 1'h0 : _GEN_825; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1082 = 6'h3a == rb_index ? 1'h0 : _GEN_826; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1083 = 6'h3b == rb_index ? 1'h0 : _GEN_827; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1084 = 6'h3c == rb_index ? 1'h0 : _GEN_828; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1085 = 6'h3d == rb_index ? 1'h0 : _GEN_829; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1086 = 6'h3e == rb_index ? 1'h0 : _GEN_830; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _GEN_1087 = 6'h3f == rb_index ? 1'h0 : _GEN_831; // @[Cache_Soc.scala 111:23 Cache_Soc.scala 111:23]
  wire  _T_8 = replace_way == 2'h2; // @[Cache_Soc.scala 112:30]
  wire  _GEN_1088 = _GEN_2439 | _GEN_832; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1089 = _GEN_2440 | _GEN_833; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1090 = _GEN_2441 | _GEN_834; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1091 = _GEN_2442 | _GEN_835; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1092 = _GEN_2443 | _GEN_836; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1093 = _GEN_2444 | _GEN_837; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1094 = _GEN_2445 | _GEN_838; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1095 = _GEN_2446 | _GEN_839; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1096 = _GEN_2447 | _GEN_840; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1097 = _GEN_2448 | _GEN_841; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1098 = _GEN_2449 | _GEN_842; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1099 = _GEN_2450 | _GEN_843; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1100 = _GEN_2451 | _GEN_844; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1101 = _GEN_2452 | _GEN_845; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1102 = _GEN_2453 | _GEN_846; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1103 = _GEN_2454 | _GEN_847; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1104 = _GEN_2455 | _GEN_848; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1105 = _GEN_2456 | _GEN_849; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1106 = _GEN_2457 | _GEN_850; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1107 = _GEN_2458 | _GEN_851; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1108 = _GEN_2459 | _GEN_852; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1109 = _GEN_2460 | _GEN_853; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1110 = _GEN_2461 | _GEN_854; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1111 = _GEN_2462 | _GEN_855; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1112 = _GEN_2463 | _GEN_856; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1113 = _GEN_2464 | _GEN_857; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1114 = _GEN_2465 | _GEN_858; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1115 = _GEN_2466 | _GEN_859; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1116 = _GEN_2467 | _GEN_860; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1117 = _GEN_2468 | _GEN_861; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1118 = _GEN_2469 | _GEN_862; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1119 = _GEN_2470 | _GEN_863; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1120 = _GEN_2471 | _GEN_864; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1121 = _GEN_2472 | _GEN_865; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1122 = _GEN_2473 | _GEN_866; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1123 = _GEN_2474 | _GEN_867; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1124 = _GEN_2475 | _GEN_868; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1125 = _GEN_2476 | _GEN_869; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1126 = _GEN_2477 | _GEN_870; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1127 = _GEN_2478 | _GEN_871; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1128 = _GEN_2479 | _GEN_872; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1129 = _GEN_2480 | _GEN_873; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1130 = _GEN_2481 | _GEN_874; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1131 = _GEN_2482 | _GEN_875; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1132 = _GEN_2483 | _GEN_876; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1133 = _GEN_2484 | _GEN_877; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1134 = _GEN_2485 | _GEN_878; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1135 = _GEN_2486 | _GEN_879; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1136 = _GEN_2487 | _GEN_880; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1137 = _GEN_2488 | _GEN_881; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1138 = _GEN_2489 | _GEN_882; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1139 = _GEN_2490 | _GEN_883; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1140 = _GEN_2491 | _GEN_884; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1141 = _GEN_2492 | _GEN_885; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1142 = _GEN_2493 | _GEN_886; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1143 = _GEN_2494 | _GEN_887; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1144 = _GEN_2495 | _GEN_888; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1145 = _GEN_2496 | _GEN_889; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1146 = _GEN_2497 | _GEN_890; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1147 = _GEN_2498 | _GEN_891; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1148 = _GEN_2499 | _GEN_892; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1149 = _GEN_2500 | _GEN_893; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1150 = _GEN_2501 | _GEN_894; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _GEN_1151 = _GEN_2502 | _GEN_895; // @[Cache_Soc.scala 113:23 Cache_Soc.scala 113:23]
  wire  _T_9 = replace_way == 2'h3; // @[Cache_Soc.scala 114:30]
  wire  _GEN_1152 = 6'h0 == rb_index ? 1'h0 : _GEN_832; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1153 = 6'h1 == rb_index ? 1'h0 : _GEN_833; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1154 = 6'h2 == rb_index ? 1'h0 : _GEN_834; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1155 = 6'h3 == rb_index ? 1'h0 : _GEN_835; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1156 = 6'h4 == rb_index ? 1'h0 : _GEN_836; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1157 = 6'h5 == rb_index ? 1'h0 : _GEN_837; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1158 = 6'h6 == rb_index ? 1'h0 : _GEN_838; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1159 = 6'h7 == rb_index ? 1'h0 : _GEN_839; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1160 = 6'h8 == rb_index ? 1'h0 : _GEN_840; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1161 = 6'h9 == rb_index ? 1'h0 : _GEN_841; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1162 = 6'ha == rb_index ? 1'h0 : _GEN_842; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1163 = 6'hb == rb_index ? 1'h0 : _GEN_843; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1164 = 6'hc == rb_index ? 1'h0 : _GEN_844; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1165 = 6'hd == rb_index ? 1'h0 : _GEN_845; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1166 = 6'he == rb_index ? 1'h0 : _GEN_846; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1167 = 6'hf == rb_index ? 1'h0 : _GEN_847; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1168 = 6'h10 == rb_index ? 1'h0 : _GEN_848; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1169 = 6'h11 == rb_index ? 1'h0 : _GEN_849; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1170 = 6'h12 == rb_index ? 1'h0 : _GEN_850; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1171 = 6'h13 == rb_index ? 1'h0 : _GEN_851; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1172 = 6'h14 == rb_index ? 1'h0 : _GEN_852; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1173 = 6'h15 == rb_index ? 1'h0 : _GEN_853; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1174 = 6'h16 == rb_index ? 1'h0 : _GEN_854; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1175 = 6'h17 == rb_index ? 1'h0 : _GEN_855; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1176 = 6'h18 == rb_index ? 1'h0 : _GEN_856; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1177 = 6'h19 == rb_index ? 1'h0 : _GEN_857; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1178 = 6'h1a == rb_index ? 1'h0 : _GEN_858; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1179 = 6'h1b == rb_index ? 1'h0 : _GEN_859; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1180 = 6'h1c == rb_index ? 1'h0 : _GEN_860; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1181 = 6'h1d == rb_index ? 1'h0 : _GEN_861; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1182 = 6'h1e == rb_index ? 1'h0 : _GEN_862; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1183 = 6'h1f == rb_index ? 1'h0 : _GEN_863; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1184 = 6'h20 == rb_index ? 1'h0 : _GEN_864; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1185 = 6'h21 == rb_index ? 1'h0 : _GEN_865; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1186 = 6'h22 == rb_index ? 1'h0 : _GEN_866; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1187 = 6'h23 == rb_index ? 1'h0 : _GEN_867; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1188 = 6'h24 == rb_index ? 1'h0 : _GEN_868; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1189 = 6'h25 == rb_index ? 1'h0 : _GEN_869; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1190 = 6'h26 == rb_index ? 1'h0 : _GEN_870; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1191 = 6'h27 == rb_index ? 1'h0 : _GEN_871; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1192 = 6'h28 == rb_index ? 1'h0 : _GEN_872; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1193 = 6'h29 == rb_index ? 1'h0 : _GEN_873; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1194 = 6'h2a == rb_index ? 1'h0 : _GEN_874; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1195 = 6'h2b == rb_index ? 1'h0 : _GEN_875; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1196 = 6'h2c == rb_index ? 1'h0 : _GEN_876; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1197 = 6'h2d == rb_index ? 1'h0 : _GEN_877; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1198 = 6'h2e == rb_index ? 1'h0 : _GEN_878; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1199 = 6'h2f == rb_index ? 1'h0 : _GEN_879; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1200 = 6'h30 == rb_index ? 1'h0 : _GEN_880; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1201 = 6'h31 == rb_index ? 1'h0 : _GEN_881; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1202 = 6'h32 == rb_index ? 1'h0 : _GEN_882; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1203 = 6'h33 == rb_index ? 1'h0 : _GEN_883; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1204 = 6'h34 == rb_index ? 1'h0 : _GEN_884; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1205 = 6'h35 == rb_index ? 1'h0 : _GEN_885; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1206 = 6'h36 == rb_index ? 1'h0 : _GEN_886; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1207 = 6'h37 == rb_index ? 1'h0 : _GEN_887; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1208 = 6'h38 == rb_index ? 1'h0 : _GEN_888; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1209 = 6'h39 == rb_index ? 1'h0 : _GEN_889; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1210 = 6'h3a == rb_index ? 1'h0 : _GEN_890; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1211 = 6'h3b == rb_index ? 1'h0 : _GEN_891; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1212 = 6'h3c == rb_index ? 1'h0 : _GEN_892; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1213 = 6'h3d == rb_index ? 1'h0 : _GEN_893; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1214 = 6'h3e == rb_index ? 1'h0 : _GEN_894; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1215 = 6'h3f == rb_index ? 1'h0 : _GEN_895; // @[Cache_Soc.scala 115:23 Cache_Soc.scala 115:23]
  wire  _GEN_1216 = replace_way == 2'h3 ? _GEN_1152 : _GEN_832; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1217 = replace_way == 2'h3 ? _GEN_1153 : _GEN_833; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1218 = replace_way == 2'h3 ? _GEN_1154 : _GEN_834; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1219 = replace_way == 2'h3 ? _GEN_1155 : _GEN_835; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1220 = replace_way == 2'h3 ? _GEN_1156 : _GEN_836; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1221 = replace_way == 2'h3 ? _GEN_1157 : _GEN_837; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1222 = replace_way == 2'h3 ? _GEN_1158 : _GEN_838; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1223 = replace_way == 2'h3 ? _GEN_1159 : _GEN_839; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1224 = replace_way == 2'h3 ? _GEN_1160 : _GEN_840; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1225 = replace_way == 2'h3 ? _GEN_1161 : _GEN_841; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1226 = replace_way == 2'h3 ? _GEN_1162 : _GEN_842; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1227 = replace_way == 2'h3 ? _GEN_1163 : _GEN_843; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1228 = replace_way == 2'h3 ? _GEN_1164 : _GEN_844; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1229 = replace_way == 2'h3 ? _GEN_1165 : _GEN_845; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1230 = replace_way == 2'h3 ? _GEN_1166 : _GEN_846; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1231 = replace_way == 2'h3 ? _GEN_1167 : _GEN_847; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1232 = replace_way == 2'h3 ? _GEN_1168 : _GEN_848; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1233 = replace_way == 2'h3 ? _GEN_1169 : _GEN_849; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1234 = replace_way == 2'h3 ? _GEN_1170 : _GEN_850; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1235 = replace_way == 2'h3 ? _GEN_1171 : _GEN_851; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1236 = replace_way == 2'h3 ? _GEN_1172 : _GEN_852; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1237 = replace_way == 2'h3 ? _GEN_1173 : _GEN_853; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1238 = replace_way == 2'h3 ? _GEN_1174 : _GEN_854; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1239 = replace_way == 2'h3 ? _GEN_1175 : _GEN_855; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1240 = replace_way == 2'h3 ? _GEN_1176 : _GEN_856; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1241 = replace_way == 2'h3 ? _GEN_1177 : _GEN_857; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1242 = replace_way == 2'h3 ? _GEN_1178 : _GEN_858; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1243 = replace_way == 2'h3 ? _GEN_1179 : _GEN_859; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1244 = replace_way == 2'h3 ? _GEN_1180 : _GEN_860; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1245 = replace_way == 2'h3 ? _GEN_1181 : _GEN_861; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1246 = replace_way == 2'h3 ? _GEN_1182 : _GEN_862; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1247 = replace_way == 2'h3 ? _GEN_1183 : _GEN_863; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1248 = replace_way == 2'h3 ? _GEN_1184 : _GEN_864; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1249 = replace_way == 2'h3 ? _GEN_1185 : _GEN_865; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1250 = replace_way == 2'h3 ? _GEN_1186 : _GEN_866; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1251 = replace_way == 2'h3 ? _GEN_1187 : _GEN_867; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1252 = replace_way == 2'h3 ? _GEN_1188 : _GEN_868; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1253 = replace_way == 2'h3 ? _GEN_1189 : _GEN_869; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1254 = replace_way == 2'h3 ? _GEN_1190 : _GEN_870; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1255 = replace_way == 2'h3 ? _GEN_1191 : _GEN_871; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1256 = replace_way == 2'h3 ? _GEN_1192 : _GEN_872; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1257 = replace_way == 2'h3 ? _GEN_1193 : _GEN_873; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1258 = replace_way == 2'h3 ? _GEN_1194 : _GEN_874; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1259 = replace_way == 2'h3 ? _GEN_1195 : _GEN_875; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1260 = replace_way == 2'h3 ? _GEN_1196 : _GEN_876; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1261 = replace_way == 2'h3 ? _GEN_1197 : _GEN_877; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1262 = replace_way == 2'h3 ? _GEN_1198 : _GEN_878; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1263 = replace_way == 2'h3 ? _GEN_1199 : _GEN_879; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1264 = replace_way == 2'h3 ? _GEN_1200 : _GEN_880; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1265 = replace_way == 2'h3 ? _GEN_1201 : _GEN_881; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1266 = replace_way == 2'h3 ? _GEN_1202 : _GEN_882; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1267 = replace_way == 2'h3 ? _GEN_1203 : _GEN_883; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1268 = replace_way == 2'h3 ? _GEN_1204 : _GEN_884; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1269 = replace_way == 2'h3 ? _GEN_1205 : _GEN_885; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1270 = replace_way == 2'h3 ? _GEN_1206 : _GEN_886; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1271 = replace_way == 2'h3 ? _GEN_1207 : _GEN_887; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1272 = replace_way == 2'h3 ? _GEN_1208 : _GEN_888; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1273 = replace_way == 2'h3 ? _GEN_1209 : _GEN_889; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1274 = replace_way == 2'h3 ? _GEN_1210 : _GEN_890; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1275 = replace_way == 2'h3 ? _GEN_1211 : _GEN_891; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1276 = replace_way == 2'h3 ? _GEN_1212 : _GEN_892; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1277 = replace_way == 2'h3 ? _GEN_1213 : _GEN_893; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1278 = replace_way == 2'h3 ? _GEN_1214 : _GEN_894; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1279 = replace_way == 2'h3 ? _GEN_1215 : _GEN_895; // @[Cache_Soc.scala 114:39]
  wire  _GEN_1280 = replace_way == 2'h2 ? _GEN_1088 : _GEN_1216; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1281 = replace_way == 2'h2 ? _GEN_1089 : _GEN_1217; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1282 = replace_way == 2'h2 ? _GEN_1090 : _GEN_1218; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1283 = replace_way == 2'h2 ? _GEN_1091 : _GEN_1219; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1284 = replace_way == 2'h2 ? _GEN_1092 : _GEN_1220; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1285 = replace_way == 2'h2 ? _GEN_1093 : _GEN_1221; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1286 = replace_way == 2'h2 ? _GEN_1094 : _GEN_1222; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1287 = replace_way == 2'h2 ? _GEN_1095 : _GEN_1223; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1288 = replace_way == 2'h2 ? _GEN_1096 : _GEN_1224; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1289 = replace_way == 2'h2 ? _GEN_1097 : _GEN_1225; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1290 = replace_way == 2'h2 ? _GEN_1098 : _GEN_1226; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1291 = replace_way == 2'h2 ? _GEN_1099 : _GEN_1227; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1292 = replace_way == 2'h2 ? _GEN_1100 : _GEN_1228; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1293 = replace_way == 2'h2 ? _GEN_1101 : _GEN_1229; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1294 = replace_way == 2'h2 ? _GEN_1102 : _GEN_1230; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1295 = replace_way == 2'h2 ? _GEN_1103 : _GEN_1231; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1296 = replace_way == 2'h2 ? _GEN_1104 : _GEN_1232; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1297 = replace_way == 2'h2 ? _GEN_1105 : _GEN_1233; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1298 = replace_way == 2'h2 ? _GEN_1106 : _GEN_1234; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1299 = replace_way == 2'h2 ? _GEN_1107 : _GEN_1235; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1300 = replace_way == 2'h2 ? _GEN_1108 : _GEN_1236; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1301 = replace_way == 2'h2 ? _GEN_1109 : _GEN_1237; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1302 = replace_way == 2'h2 ? _GEN_1110 : _GEN_1238; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1303 = replace_way == 2'h2 ? _GEN_1111 : _GEN_1239; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1304 = replace_way == 2'h2 ? _GEN_1112 : _GEN_1240; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1305 = replace_way == 2'h2 ? _GEN_1113 : _GEN_1241; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1306 = replace_way == 2'h2 ? _GEN_1114 : _GEN_1242; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1307 = replace_way == 2'h2 ? _GEN_1115 : _GEN_1243; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1308 = replace_way == 2'h2 ? _GEN_1116 : _GEN_1244; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1309 = replace_way == 2'h2 ? _GEN_1117 : _GEN_1245; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1310 = replace_way == 2'h2 ? _GEN_1118 : _GEN_1246; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1311 = replace_way == 2'h2 ? _GEN_1119 : _GEN_1247; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1312 = replace_way == 2'h2 ? _GEN_1120 : _GEN_1248; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1313 = replace_way == 2'h2 ? _GEN_1121 : _GEN_1249; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1314 = replace_way == 2'h2 ? _GEN_1122 : _GEN_1250; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1315 = replace_way == 2'h2 ? _GEN_1123 : _GEN_1251; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1316 = replace_way == 2'h2 ? _GEN_1124 : _GEN_1252; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1317 = replace_way == 2'h2 ? _GEN_1125 : _GEN_1253; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1318 = replace_way == 2'h2 ? _GEN_1126 : _GEN_1254; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1319 = replace_way == 2'h2 ? _GEN_1127 : _GEN_1255; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1320 = replace_way == 2'h2 ? _GEN_1128 : _GEN_1256; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1321 = replace_way == 2'h2 ? _GEN_1129 : _GEN_1257; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1322 = replace_way == 2'h2 ? _GEN_1130 : _GEN_1258; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1323 = replace_way == 2'h2 ? _GEN_1131 : _GEN_1259; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1324 = replace_way == 2'h2 ? _GEN_1132 : _GEN_1260; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1325 = replace_way == 2'h2 ? _GEN_1133 : _GEN_1261; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1326 = replace_way == 2'h2 ? _GEN_1134 : _GEN_1262; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1327 = replace_way == 2'h2 ? _GEN_1135 : _GEN_1263; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1328 = replace_way == 2'h2 ? _GEN_1136 : _GEN_1264; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1329 = replace_way == 2'h2 ? _GEN_1137 : _GEN_1265; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1330 = replace_way == 2'h2 ? _GEN_1138 : _GEN_1266; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1331 = replace_way == 2'h2 ? _GEN_1139 : _GEN_1267; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1332 = replace_way == 2'h2 ? _GEN_1140 : _GEN_1268; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1333 = replace_way == 2'h2 ? _GEN_1141 : _GEN_1269; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1334 = replace_way == 2'h2 ? _GEN_1142 : _GEN_1270; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1335 = replace_way == 2'h2 ? _GEN_1143 : _GEN_1271; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1336 = replace_way == 2'h2 ? _GEN_1144 : _GEN_1272; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1337 = replace_way == 2'h2 ? _GEN_1145 : _GEN_1273; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1338 = replace_way == 2'h2 ? _GEN_1146 : _GEN_1274; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1339 = replace_way == 2'h2 ? _GEN_1147 : _GEN_1275; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1340 = replace_way == 2'h2 ? _GEN_1148 : _GEN_1276; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1341 = replace_way == 2'h2 ? _GEN_1149 : _GEN_1277; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1342 = replace_way == 2'h2 ? _GEN_1150 : _GEN_1278; // @[Cache_Soc.scala 112:39]
  wire  _GEN_1343 = replace_way == 2'h2 ? _GEN_1151 : _GEN_1279; // @[Cache_Soc.scala 112:39]
  wire  _addr_ok_T = state == 3'h0; // @[Cache_Soc.scala 156:22]
  wire  conflict = wb_state & io_in_valid; // @[Cache_Soc.scala 155:38]
  wire  addr_ok = (state == 3'h0 | _T_1) & io_in_valid & ~conflict; // @[Cache_Soc.scala 156:80]
  wire  _T_10 = io_in_valid & addr_ok; // @[Cache_Soc.scala 127:18]
  wire  _T_14 = _T_1 & rb_op; // @[Cache_Soc.scala 138:41]
  wire [3:0] _wb_hitway_T = {hit_3,hit_2,hit_1,hit_0}; // @[OneHot.scala 22:45]
  wire [1:0] wb_hitway_hi_1 = _wb_hitway_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] wb_hitway_lo_1 = _wb_hitway_T[1:0]; // @[OneHot.scala 31:18]
  wire  wb_hitway_hi_2 = |wb_hitway_hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _wb_hitway_T_1 = wb_hitway_hi_1 | wb_hitway_lo_1; // @[OneHot.scala 32:28]
  wire  wb_hitway_lo_2 = _wb_hitway_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] _wb_hitway_T_2 = {wb_hitway_hi_2,wb_hitway_lo_2}; // @[Cat.scala 30:58]
  wire  _GEN_1998 = 2'h1 == replace_way ? valid_1 : valid_0; // @[Cache_Soc.scala 149:19 Cache_Soc.scala 149:19]
  wire  dirty_0 = meta_0_io_dirty_r;
  wire  dirty_1 = meta_1_io_dirty_r;
  wire  _GEN_2002 = 2'h1 == replace_way ? dirty_1 : dirty_0; // @[Cache_Soc.scala 150:19 Cache_Soc.scala 150:19]
  wire  dirty_2 = meta_2_io_dirty_r;
  wire  dirty_3 = meta_3_io_dirty_r;
  wire [21:0] _GEN_2006 = 2'h1 == replace_way ? tag_1 : tag_0; // @[Cache_Soc.scala 151:17 Cache_Soc.scala 151:17]
  wire [127:0] _GEN_2010 = 2'h1 == replace_way ? io_sram_1_rdata : io_sram_0_rdata; // @[Cache_Soc.scala 152:18 Cache_Soc.scala 152:18]
  wire  _io_in_data_ok_T_4 = rb_uncache & rb_op; // @[Cache_Soc.scala 157:90]
  wire  _io_in_data_ok_T_6 = rb_uncache & rb_op & io_out_wr_ok | io_out_ret_valid; // @[Cache_Soc.scala 157:123]
  wire [63:0] _load_res_T_3 = rb_offset[3] ? io_sram_0_rdata[127:64] : io_sram_0_rdata[63:0]; // @[Cache_Soc.scala 162:22]
  wire [63:0] _GEN_2017 = hit_0 ? _load_res_T_3 : 64'h0; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 162:16]
  wire [127:0] _GEN_2018 = hit_0 ? io_sram_0_rdata : 128'h0; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 163:17]
  wire [63:0] _load_res_T_7 = rb_offset[3] ? io_sram_1_rdata[127:64] : io_sram_1_rdata[63:0]; // @[Cache_Soc.scala 162:22]
  wire [63:0] _GEN_2019 = hit_1 ? _load_res_T_7 : _GEN_2017; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 162:16]
  wire [127:0] _GEN_2020 = hit_1 ? io_sram_1_rdata : _GEN_2018; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 163:17]
  wire [63:0] _load_res_T_11 = rb_offset[3] ? io_sram_2_rdata[127:64] : io_sram_2_rdata[63:0]; // @[Cache_Soc.scala 162:22]
  wire [63:0] _GEN_2021 = hit_2 ? _load_res_T_11 : _GEN_2019; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 162:16]
  wire [127:0] _GEN_2022 = hit_2 ? io_sram_2_rdata : _GEN_2020; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 163:17]
  wire [63:0] _load_res_T_15 = rb_offset[3] ? io_sram_3_rdata[127:64] : io_sram_3_rdata[63:0]; // @[Cache_Soc.scala 162:22]
  wire [63:0] load_res = hit_3 ? _load_res_T_15 : _GEN_2021; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 162:16]
  wire [127:0] load_inst = hit_3 ? io_sram_3_rdata : _GEN_2022; // @[Cache_Soc.scala 161:19 Cache_Soc.scala 163:17]
  wire [63:0] rd_rdata = rb_offset[3] | rb_uncache ? io_out_ret_data[127:64] : io_out_ret_data[63:0]; // @[Cache_Soc.scala 168:18]
  wire [127:0] _rd_inst_T = {io_out_ret_data[127:64],io_out_ret_data[127:64]}; // @[Cat.scala 30:58]
  wire [127:0] rd_inst = rb_uncache ? _rd_inst_T : io_out_ret_data; // @[Cache_Soc.scala 169:17]
  wire [63:0] _io_in_rdata_T_4 = _T_3 ? rd_rdata : 64'h0; // @[Cache_Soc.scala 170:65]
  wire [127:0] _io_in_inst_T_4 = _T_3 ? rd_inst : 128'h0; // @[Cache_Soc.scala 171:65]
  wire [2:0] _io_out_wr_size_T = rb_uncache ? 3'h2 : 3'h3; // @[Cache_Soc.scala 176:21]
  wire [31:0] _io_out_wr_addr_T = {rb_tag,rb_index,rb_offset}; // @[Cat.scala 30:58]
  wire [31:0] _io_out_wr_addr_T_1 = {replace_tag,rb_index,4'h0}; // @[Cat.scala 30:58]
  wire [31:0] _io_out_wr_addr_T_2 = rb_uncache ? _io_out_wr_addr_T : _io_out_wr_addr_T_1; // @[Cache_Soc.scala 177:21]
  wire [7:0] _io_out_wr_wstrb_T = rb_uncache ? rb_wstrb : 8'hff; // @[Cache_Soc.scala 178:22]
  wire [127:0] _io_out_wr_data_T = {rb_wdata,rb_wdata}; // @[Cat.scala 30:58]
  wire [127:0] _io_out_wr_data_T_1 = rb_uncache ? _io_out_wr_data_T : replace_data; // @[Cache_Soc.scala 179:21]
  wire [31:0] _io_out_rd_addr_T_1 = {rb_tag,rb_index,4'h0}; // @[Cat.scala 30:58]
  wire  _T_18 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_20 = ~in_uncache; // @[Cache_Soc.scala 188:15]
  wire [5:0] _GEN_2026 = ~in_uncache ? in_index : 6'h0; // @[Cache_Soc.scala 188:28 Cache_Soc.scala 191:26 Cache_Soc.scala 19:12]
  wire  _GEN_2028 = _T_10 & _T_20; // @[Cache_Soc.scala 186:34 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2029 = _T_10 ? _GEN_2026 : 6'h0; // @[Cache_Soc.scala 186:34 Cache_Soc.scala 19:12]
  wire  _T_21 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_2032 = cache_hit ? 3'h0 : 3'h2; // @[Cache_Soc.scala 207:31 Cache_Soc.scala 208:15 Cache_Soc.scala 210:15]
  wire  _GEN_2034 = cache_hit & _T_10 & _T_20; // @[Cache_Soc.scala 198:49 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2035 = cache_hit & _T_10 ? _GEN_2026 : 6'h0; // @[Cache_Soc.scala 198:49 Cache_Soc.scala 19:12]
  wire  _T_25 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_33 = io_out_wr_req & io_out_wr_rdy; // @[Cache_Soc.scala 218:31]
  wire [2:0] _GEN_2036 = io_out_wr_req & io_out_wr_rdy ? 3'h3 : state; // @[Cache_Soc.scala 218:46 Cache_Soc.scala 219:15 Cache_Soc.scala 41:22]
  wire [2:0] _GEN_2037 = _cache_hit_T_2 & ~(replace_valid & replace_dirty) | rb_uncache & ~rb_op ? 3'h3 : _GEN_2036; // @[Cache_Soc.scala 215:101 Cache_Soc.scala 216:15]
  wire  _GEN_2038 = _cache_hit_T_2 & ~(replace_valid & replace_dirty) | rb_uncache & ~rb_op ? 1'h0 : 1'h1; // @[Cache_Soc.scala 215:101 Cache_Soc.scala 217:20 Cache_Soc.scala 214:18]
  wire  _T_34 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_2039 = io_out_rd_req & io_out_rd_rdy ? 3'h4 : state; // @[Cache_Soc.scala 227:46 Cache_Soc.scala 228:15 Cache_Soc.scala 41:22]
  wire [2:0] _GEN_2040 = _io_in_data_ok_T_4 ? 3'h4 : _GEN_2039; // @[Cache_Soc.scala 224:46 Cache_Soc.scala 225:15]
  wire  _GEN_2041 = _io_in_data_ok_T_4 ? 1'h0 : 1'h1; // @[Cache_Soc.scala 224:46 Cache_Soc.scala 226:20 Cache_Soc.scala 223:18]
  wire  _T_38 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_2042 = _io_in_data_ok_T_6 ? 3'h0 : state; // @[Cache_Soc.scala 238:74 Cache_Soc.scala 239:15 Cache_Soc.scala 41:22]
  wire  _T_46 = _plru0_T_1 & io_out_ret_valid & _cache_hit_T_2; // @[Cache_Soc.scala 243:52]
  wire [7:0] io_sram_0_wdata_lo_lo_lo = rb_wstrb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_lo_lo_hi = rb_wstrb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_lo_hi_lo = rb_wstrb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_lo_hi_hi = rb_wstrb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_lo_lo = rb_wstrb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_lo_hi = rb_wstrb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_hi_lo = rb_wstrb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_hi_hi = rb_wstrb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_sram_0_wdata_T_18 = {io_sram_0_wdata_hi_hi_hi,io_sram_0_wdata_hi_hi_lo,io_sram_0_wdata_hi_lo_hi,
    io_sram_0_wdata_hi_lo_lo,io_sram_0_wdata_lo_hi_hi,io_sram_0_wdata_lo_hi_lo,io_sram_0_wdata_lo_lo_hi,
    io_sram_0_wdata_lo_lo_lo}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_0_wdata_T_19 = rb_wdata & _io_sram_0_wdata_T_18; // @[MAP.scala 10:14]
  wire [63:0] _io_sram_0_wdata_T_20 = ~_io_sram_0_wdata_T_18; // @[MAP.scala 10:35]
  wire [63:0] _io_sram_0_wdata_T_21 = io_out_ret_data[127:64] & _io_sram_0_wdata_T_20; // @[MAP.scala 10:33]
  wire [63:0] io_sram_0_wdata_hi_1 = _io_sram_0_wdata_T_19 | _io_sram_0_wdata_T_21; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_0_wdata_T_22 = {io_sram_0_wdata_hi_1,io_out_ret_data[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_0_wdata_T_43 = io_out_ret_data[63:0] & _io_sram_0_wdata_T_20; // @[MAP.scala 10:33]
  wire [63:0] io_sram_0_wdata_lo_3 = _io_sram_0_wdata_T_19 | _io_sram_0_wdata_T_43; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_0_wdata_T_44 = {io_out_ret_data[127:64],io_sram_0_wdata_lo_3}; // @[Cat.scala 30:58]
  wire [127:0] _io_sram_0_wdata_T_45 = rb_offset[3] ? _io_sram_0_wdata_T_22 : _io_sram_0_wdata_T_44; // @[Cache_Soc.scala 248:33]
  wire [127:0] _GEN_2043 = rb_op ? _io_sram_0_wdata_T_45 : io_out_ret_data; // @[Cache_Soc.scala 247:34 Cache_Soc.scala 248:27 Cache_Soc.scala 252:27]
  wire [5:0] _GEN_2045 = _plru0_T_1 & io_out_ret_valid & _cache_hit_T_2 ? rb_index : 6'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 246:24 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2046 = _plru0_T_1 & io_out_ret_valid & _cache_hit_T_2 ? _GEN_2043 : 128'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2047 = _plru0_T_1 & io_out_ret_valid & _cache_hit_T_2 ? rb_tag : 22'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 255:28 Cache_Soc.scala 30:16]
  wire  _GEN_2048 = _plru0_T_1 & io_out_ret_valid & _cache_hit_T_2 & rb_op; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 258:30 Cache_Soc.scala 32:18]
  wire  _T_51 = _plru0_T_2 & io_out_ret_valid & _cache_hit_T_2; // @[Cache_Soc.scala 243:52]
  wire [5:0] _GEN_2051 = _plru0_T_2 & io_out_ret_valid & _cache_hit_T_2 ? rb_index : 6'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 246:24 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2052 = _plru0_T_2 & io_out_ret_valid & _cache_hit_T_2 ? _GEN_2043 : 128'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2053 = _plru0_T_2 & io_out_ret_valid & _cache_hit_T_2 ? rb_tag : 22'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 255:28 Cache_Soc.scala 30:16]
  wire  _GEN_2054 = _plru0_T_2 & io_out_ret_valid & _cache_hit_T_2 & rb_op; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 258:30 Cache_Soc.scala 32:18]
  wire  _T_56 = _T_8 & io_out_ret_valid & _cache_hit_T_2; // @[Cache_Soc.scala 243:52]
  wire [5:0] _GEN_2057 = _T_8 & io_out_ret_valid & _cache_hit_T_2 ? rb_index : 6'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 246:24 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2058 = _T_8 & io_out_ret_valid & _cache_hit_T_2 ? _GEN_2043 : 128'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2059 = _T_8 & io_out_ret_valid & _cache_hit_T_2 ? rb_tag : 22'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 255:28 Cache_Soc.scala 30:16]
  wire  _GEN_2060 = _T_8 & io_out_ret_valid & _cache_hit_T_2 & rb_op; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 258:30 Cache_Soc.scala 32:18]
  wire  _T_61 = _T_9 & io_out_ret_valid & _cache_hit_T_2; // @[Cache_Soc.scala 243:52]
  wire [5:0] _GEN_2063 = _T_9 & io_out_ret_valid & _cache_hit_T_2 ? rb_index : 6'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 246:24 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2064 = _T_9 & io_out_ret_valid & _cache_hit_T_2 ? _GEN_2043 : 128'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2065 = _T_9 & io_out_ret_valid & _cache_hit_T_2 ? rb_tag : 22'h0; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 255:28 Cache_Soc.scala 30:16]
  wire  _GEN_2066 = _T_9 & io_out_ret_valid & _cache_hit_T_2 & rb_op; // @[Cache_Soc.scala 243:68 Cache_Soc.scala 258:30 Cache_Soc.scala 32:18]
  wire [2:0] _GEN_2067 = _T_38 ? _GEN_2042 : state; // @[Conditional.scala 39:67 Cache_Soc.scala 41:22]
  wire [5:0] _GEN_2069 = _T_38 ? _GEN_2045 : 6'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2070 = _T_38 ? _GEN_2046 : 128'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2071 = _T_38 ? _GEN_2047 : 22'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire [5:0] _GEN_2074 = _T_38 ? _GEN_2051 : 6'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2075 = _T_38 ? _GEN_2052 : 128'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2076 = _T_38 ? _GEN_2053 : 22'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire [5:0] _GEN_2079 = _T_38 ? _GEN_2057 : 6'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2080 = _T_38 ? _GEN_2058 : 128'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2081 = _T_38 ? _GEN_2059 : 22'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire [5:0] _GEN_2084 = _T_38 ? _GEN_2063 : 6'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2085 = _T_38 ? _GEN_2064 : 128'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2086 = _T_38 ? _GEN_2065 : 22'h0; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire [2:0] _GEN_2089 = _T_34 ? _GEN_2040 : _GEN_2067; // @[Conditional.scala 39:67]
  wire  _GEN_2090 = _T_34 ? 1'h0 : _T_38 & _T_46; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2091 = _T_34 ? 6'h0 : _GEN_2069; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2092 = _T_34 ? 128'h0 : _GEN_2070; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2093 = _T_34 ? 22'h0 : _GEN_2071; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2094 = _T_34 ? 1'h0 : _T_38 & _GEN_2048; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2095 = _T_34 ? 1'h0 : _T_38 & _T_51; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2096 = _T_34 ? 6'h0 : _GEN_2074; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2097 = _T_34 ? 128'h0 : _GEN_2075; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2098 = _T_34 ? 22'h0 : _GEN_2076; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2099 = _T_34 ? 1'h0 : _T_38 & _GEN_2054; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2100 = _T_34 ? 1'h0 : _T_38 & _T_56; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2101 = _T_34 ? 6'h0 : _GEN_2079; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2102 = _T_34 ? 128'h0 : _GEN_2080; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2103 = _T_34 ? 22'h0 : _GEN_2081; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2104 = _T_34 ? 1'h0 : _T_38 & _GEN_2060; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2105 = _T_34 ? 1'h0 : _T_38 & _T_61; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2106 = _T_34 ? 6'h0 : _GEN_2084; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2107 = _T_34 ? 128'h0 : _GEN_2085; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2108 = _T_34 ? 22'h0 : _GEN_2086; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2109 = _T_34 ? 1'h0 : _T_38 & _GEN_2066; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2112 = _T_25 ? 1'h0 : _T_34 & _GEN_2041; // @[Conditional.scala 39:67 Cache_Soc.scala 174:14]
  wire  _GEN_2113 = _T_25 ? 1'h0 : _GEN_2090; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2114 = _T_25 ? 6'h0 : _GEN_2091; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2115 = _T_25 ? 128'h0 : _GEN_2092; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2116 = _T_25 ? 22'h0 : _GEN_2093; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2117 = _T_25 ? 1'h0 : _GEN_2094; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2118 = _T_25 ? 1'h0 : _GEN_2095; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2119 = _T_25 ? 6'h0 : _GEN_2096; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2120 = _T_25 ? 128'h0 : _GEN_2097; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2121 = _T_25 ? 22'h0 : _GEN_2098; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2122 = _T_25 ? 1'h0 : _GEN_2099; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2123 = _T_25 ? 1'h0 : _GEN_2100; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2124 = _T_25 ? 6'h0 : _GEN_2101; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2125 = _T_25 ? 128'h0 : _GEN_2102; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2126 = _T_25 ? 22'h0 : _GEN_2103; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2127 = _T_25 ? 1'h0 : _GEN_2104; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2128 = _T_25 ? 1'h0 : _GEN_2105; // @[Conditional.scala 39:67 Cache_Soc.scala 17:10]
  wire [5:0] _GEN_2129 = _T_25 ? 6'h0 : _GEN_2106; // @[Conditional.scala 39:67 Cache_Soc.scala 19:12]
  wire [127:0] _GEN_2130 = _T_25 ? 128'h0 : _GEN_2107; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2131 = _T_25 ? 22'h0 : _GEN_2108; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2132 = _T_25 ? 1'h0 : _GEN_2109; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2134 = _T_21 ? _GEN_2034 : _GEN_2113; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2135 = _T_21 ? _GEN_2035 : _GEN_2114; // @[Conditional.scala 39:67]
  wire  _GEN_2136 = _T_21 ? _GEN_2034 : _GEN_2118; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2137 = _T_21 ? _GEN_2035 : _GEN_2119; // @[Conditional.scala 39:67]
  wire  _GEN_2138 = _T_21 ? _GEN_2034 : _GEN_2123; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2139 = _T_21 ? _GEN_2035 : _GEN_2124; // @[Conditional.scala 39:67]
  wire  _GEN_2140 = _T_21 ? _GEN_2034 : _GEN_2128; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2141 = _T_21 ? _GEN_2035 : _GEN_2129; // @[Conditional.scala 39:67]
  wire  _GEN_2142 = _T_21 ? 1'h0 : _T_25 & _GEN_2038; // @[Conditional.scala 39:67 Cache_Soc.scala 173:14]
  wire  _GEN_2143 = _T_21 ? 1'h0 : _GEN_2112; // @[Conditional.scala 39:67 Cache_Soc.scala 174:14]
  wire  _GEN_2144 = _T_21 ? 1'h0 : _GEN_2113; // @[Conditional.scala 39:67 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2145 = _T_21 ? 128'h0 : _GEN_2115; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2146 = _T_21 ? 22'h0 : _GEN_2116; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2147 = _T_21 ? 1'h0 : _GEN_2117; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2148 = _T_21 ? 1'h0 : _GEN_2118; // @[Conditional.scala 39:67 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2149 = _T_21 ? 128'h0 : _GEN_2120; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2150 = _T_21 ? 22'h0 : _GEN_2121; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2151 = _T_21 ? 1'h0 : _GEN_2122; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2152 = _T_21 ? 1'h0 : _GEN_2123; // @[Conditional.scala 39:67 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2153 = _T_21 ? 128'h0 : _GEN_2125; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2154 = _T_21 ? 22'h0 : _GEN_2126; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2155 = _T_21 ? 1'h0 : _GEN_2127; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2156 = _T_21 ? 1'h0 : _GEN_2128; // @[Conditional.scala 39:67 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2157 = _T_21 ? 128'h0 : _GEN_2130; // @[Conditional.scala 39:67 Cache_Soc.scala 20:13]
  wire [21:0] _GEN_2158 = _T_21 ? 22'h0 : _GEN_2131; // @[Conditional.scala 39:67 Cache_Soc.scala 30:16]
  wire  _GEN_2159 = _T_21 ? 1'h0 : _GEN_2132; // @[Conditional.scala 39:67 Cache_Soc.scala 32:18]
  wire  _GEN_2161 = _T_18 ? _GEN_2028 : _GEN_2134; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2162 = _T_18 ? _GEN_2029 : _GEN_2135; // @[Conditional.scala 40:58]
  wire  _GEN_2163 = _T_18 ? _GEN_2028 : _GEN_2136; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2164 = _T_18 ? _GEN_2029 : _GEN_2137; // @[Conditional.scala 40:58]
  wire  _GEN_2165 = _T_18 ? _GEN_2028 : _GEN_2138; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2166 = _T_18 ? _GEN_2029 : _GEN_2139; // @[Conditional.scala 40:58]
  wire  _GEN_2167 = _T_18 ? _GEN_2028 : _GEN_2140; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2168 = _T_18 ? _GEN_2029 : _GEN_2141; // @[Conditional.scala 40:58]
  wire  _GEN_2169 = _T_18 ? 1'h0 : _GEN_2142; // @[Conditional.scala 40:58 Cache_Soc.scala 173:14]
  wire  _GEN_2171 = _T_18 ? 1'h0 : _GEN_2144; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2172 = _T_18 ? 128'h0 : _GEN_2145; // @[Conditional.scala 40:58 Cache_Soc.scala 20:13]
  wire  _GEN_2174 = _T_18 ? 1'h0 : _GEN_2147; // @[Conditional.scala 40:58 Cache_Soc.scala 32:18]
  wire  _GEN_2175 = _T_18 ? 1'h0 : _GEN_2148; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2176 = _T_18 ? 128'h0 : _GEN_2149; // @[Conditional.scala 40:58 Cache_Soc.scala 20:13]
  wire  _GEN_2178 = _T_18 ? 1'h0 : _GEN_2151; // @[Conditional.scala 40:58 Cache_Soc.scala 32:18]
  wire  _GEN_2179 = _T_18 ? 1'h0 : _GEN_2152; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2180 = _T_18 ? 128'h0 : _GEN_2153; // @[Conditional.scala 40:58 Cache_Soc.scala 20:13]
  wire  _GEN_2182 = _T_18 ? 1'h0 : _GEN_2155; // @[Conditional.scala 40:58 Cache_Soc.scala 32:18]
  wire  _GEN_2183 = _T_18 ? 1'h0 : _GEN_2156; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  wire [127:0] _GEN_2184 = _T_18 ? 128'h0 : _GEN_2157; // @[Conditional.scala 40:58 Cache_Soc.scala 20:13]
  wire  _GEN_2186 = _T_18 ? 1'h0 : _GEN_2159; // @[Conditional.scala 40:58 Cache_Soc.scala 32:18]
  wire  _T_63 = ~wb_state; // @[Conditional.scala 37:30]
  wire  _GEN_2187 = hit_0 | _GEN_2161; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 271:24]
  wire [5:0] _GEN_2188 = hit_0 ? rb_index : _GEN_2162; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 272:26]
  wire  _GEN_2189 = hit_1 | _GEN_2163; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 271:24]
  wire [5:0] _GEN_2190 = hit_1 ? rb_index : _GEN_2164; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 272:26]
  wire  _GEN_2191 = hit_2 | _GEN_2165; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 271:24]
  wire [5:0] _GEN_2192 = hit_2 ? rb_index : _GEN_2166; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 272:26]
  wire  _GEN_2193 = hit_3 | _GEN_2167; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 271:24]
  wire [5:0] _GEN_2194 = hit_3 ? rb_index : _GEN_2168; // @[Cache_Soc.scala 270:25 Cache_Soc.scala 272:26]
  wire  _GEN_2195 = _T_14 | wb_state; // @[Cache_Soc.scala 267:67 Cache_Soc.scala 268:18 Cache_Soc.scala 42:25]
  wire  _GEN_2196 = _T_14 ? _GEN_2187 : _GEN_2161; // @[Cache_Soc.scala 267:67]
  wire [5:0] _GEN_2197 = _T_14 ? _GEN_2188 : _GEN_2162; // @[Cache_Soc.scala 267:67]
  wire  _GEN_2198 = _T_14 ? _GEN_2189 : _GEN_2163; // @[Cache_Soc.scala 267:67]
  wire [5:0] _GEN_2199 = _T_14 ? _GEN_2190 : _GEN_2164; // @[Cache_Soc.scala 267:67]
  wire  _GEN_2200 = _T_14 ? _GEN_2191 : _GEN_2165; // @[Cache_Soc.scala 267:67]
  wire [5:0] _GEN_2201 = _T_14 ? _GEN_2192 : _GEN_2166; // @[Cache_Soc.scala 267:67]
  wire  _GEN_2202 = _T_14 ? _GEN_2193 : _GEN_2167; // @[Cache_Soc.scala 267:67]
  wire [5:0] _GEN_2203 = _T_14 ? _GEN_2194 : _GEN_2168; // @[Cache_Soc.scala 267:67]
  wire [7:0] io_sram_0_wdata_lo_lo_lo_2 = wb_wstrb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_lo_lo_hi_2 = wb_wstrb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_lo_hi_lo_2 = wb_wstrb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_lo_hi_hi_2 = wb_wstrb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_lo_lo_2 = wb_wstrb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_lo_hi_2 = wb_wstrb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_hi_lo_2 = wb_wstrb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] io_sram_0_wdata_hi_hi_hi_2 = wb_wstrb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _io_sram_0_wdata_T_64 = {io_sram_0_wdata_hi_hi_hi_2,io_sram_0_wdata_hi_hi_lo_2,io_sram_0_wdata_hi_lo_hi_2,
    io_sram_0_wdata_hi_lo_lo_2,io_sram_0_wdata_lo_hi_hi_2,io_sram_0_wdata_lo_hi_lo_2,io_sram_0_wdata_lo_lo_hi_2,
    io_sram_0_wdata_lo_lo_lo_2}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_0_wdata_T_65 = wb_wdata & _io_sram_0_wdata_T_64; // @[MAP.scala 10:14]
  wire [63:0] _io_sram_0_wdata_T_66 = ~_io_sram_0_wdata_T_64; // @[MAP.scala 10:35]
  wire [63:0] _io_sram_0_wdata_T_67 = io_sram_0_rdata[127:64] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_0_wdata_hi_5 = _io_sram_0_wdata_T_65 | _io_sram_0_wdata_T_67; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_0_wdata_T_68 = {io_sram_0_wdata_hi_5,io_sram_0_rdata[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_0_wdata_T_89 = io_sram_0_rdata[63:0] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_0_wdata_lo_7 = _io_sram_0_wdata_T_65 | _io_sram_0_wdata_T_89; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_0_wdata_T_90 = {io_sram_0_rdata[127:64],io_sram_0_wdata_lo_7}; // @[Cat.scala 30:58]
  wire [127:0] _io_sram_0_wdata_T_91 = wb_offset[3] ? _io_sram_0_wdata_T_68 : _io_sram_0_wdata_T_90; // @[Cache_Soc.scala 284:31]
  wire  _GEN_2204 = wb_hitway == 2'h0 | _GEN_2161; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 281:22]
  wire  _GEN_2205 = wb_hitway == 2'h0 | _GEN_2171; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 282:23]
  wire [5:0] _GEN_2206 = wb_hitway == 2'h0 ? wb_index : _GEN_2162; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 283:24]
  wire [127:0] _GEN_2207 = wb_hitway == 2'h0 ? _io_sram_0_wdata_T_91 : _GEN_2172; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 284:25]
  wire  _GEN_2208 = wb_hitway == 2'h0 | _GEN_2174; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 289:30]
  wire [63:0] _io_sram_1_wdata_T_67 = io_sram_1_rdata[127:64] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_1_wdata_hi_5 = _io_sram_0_wdata_T_65 | _io_sram_1_wdata_T_67; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_1_wdata_T_68 = {io_sram_1_wdata_hi_5,io_sram_1_rdata[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_1_wdata_T_89 = io_sram_1_rdata[63:0] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_1_wdata_lo_7 = _io_sram_0_wdata_T_65 | _io_sram_1_wdata_T_89; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_1_wdata_T_90 = {io_sram_1_rdata[127:64],io_sram_1_wdata_lo_7}; // @[Cat.scala 30:58]
  wire [127:0] _io_sram_1_wdata_T_91 = wb_offset[3] ? _io_sram_1_wdata_T_68 : _io_sram_1_wdata_T_90; // @[Cache_Soc.scala 284:31]
  wire  _GEN_2209 = wb_hitway == 2'h1 | _GEN_2163; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 281:22]
  wire  _GEN_2210 = wb_hitway == 2'h1 | _GEN_2175; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 282:23]
  wire [5:0] _GEN_2211 = wb_hitway == 2'h1 ? wb_index : _GEN_2164; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 283:24]
  wire [127:0] _GEN_2212 = wb_hitway == 2'h1 ? _io_sram_1_wdata_T_91 : _GEN_2176; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 284:25]
  wire  _GEN_2213 = wb_hitway == 2'h1 | _GEN_2178; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 289:30]
  wire [63:0] _io_sram_2_wdata_T_67 = io_sram_2_rdata[127:64] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_2_wdata_hi_5 = _io_sram_0_wdata_T_65 | _io_sram_2_wdata_T_67; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_2_wdata_T_68 = {io_sram_2_wdata_hi_5,io_sram_2_rdata[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_2_wdata_T_89 = io_sram_2_rdata[63:0] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_2_wdata_lo_7 = _io_sram_0_wdata_T_65 | _io_sram_2_wdata_T_89; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_2_wdata_T_90 = {io_sram_2_rdata[127:64],io_sram_2_wdata_lo_7}; // @[Cat.scala 30:58]
  wire [127:0] _io_sram_2_wdata_T_91 = wb_offset[3] ? _io_sram_2_wdata_T_68 : _io_sram_2_wdata_T_90; // @[Cache_Soc.scala 284:31]
  wire  _GEN_2214 = wb_hitway == 2'h2 | _GEN_2165; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 281:22]
  wire  _GEN_2215 = wb_hitway == 2'h2 | _GEN_2179; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 282:23]
  wire [5:0] _GEN_2216 = wb_hitway == 2'h2 ? wb_index : _GEN_2166; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 283:24]
  wire [127:0] _GEN_2217 = wb_hitway == 2'h2 ? _io_sram_2_wdata_T_91 : _GEN_2180; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 284:25]
  wire  _GEN_2218 = wb_hitway == 2'h2 | _GEN_2182; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 289:30]
  wire [63:0] _io_sram_3_wdata_T_67 = io_sram_3_rdata[127:64] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_3_wdata_hi_5 = _io_sram_0_wdata_T_65 | _io_sram_3_wdata_T_67; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_3_wdata_T_68 = {io_sram_3_wdata_hi_5,io_sram_3_rdata[63:0]}; // @[Cat.scala 30:58]
  wire [63:0] _io_sram_3_wdata_T_89 = io_sram_3_rdata[63:0] & _io_sram_0_wdata_T_66; // @[MAP.scala 10:33]
  wire [63:0] io_sram_3_wdata_lo_7 = _io_sram_0_wdata_T_65 | _io_sram_3_wdata_T_89; // @[MAP.scala 10:22]
  wire [127:0] _io_sram_3_wdata_T_90 = {io_sram_3_rdata[127:64],io_sram_3_wdata_lo_7}; // @[Cat.scala 30:58]
  wire [127:0] _io_sram_3_wdata_T_91 = wb_offset[3] ? _io_sram_3_wdata_T_68 : _io_sram_3_wdata_T_90; // @[Cache_Soc.scala 284:31]
  wire  _GEN_2219 = wb_hitway == 2'h3 | _GEN_2167; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 281:22]
  wire  _GEN_2220 = wb_hitway == 2'h3 | _GEN_2183; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 282:23]
  wire [5:0] _GEN_2221 = wb_hitway == 2'h3 ? wb_index : _GEN_2168; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 283:24]
  wire [127:0] _GEN_2222 = wb_hitway == 2'h3 ? _io_sram_3_wdata_T_91 : _GEN_2184; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 284:25]
  wire  _GEN_2223 = wb_hitway == 2'h3 | _GEN_2186; // @[Cache_Soc.scala 280:34 Cache_Soc.scala 289:30]
  wire  _GEN_2225 = wb_state ? _GEN_2204 : _GEN_2161; // @[Conditional.scala 39:67]
  wire  _GEN_2226 = wb_state ? _GEN_2205 : _GEN_2171; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2227 = wb_state ? _GEN_2206 : _GEN_2162; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2228 = wb_state ? _GEN_2207 : _GEN_2172; // @[Conditional.scala 39:67]
  wire  _GEN_2229 = wb_state ? _GEN_2208 : _GEN_2174; // @[Conditional.scala 39:67]
  wire  _GEN_2230 = wb_state ? _GEN_2209 : _GEN_2163; // @[Conditional.scala 39:67]
  wire  _GEN_2231 = wb_state ? _GEN_2210 : _GEN_2175; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2232 = wb_state ? _GEN_2211 : _GEN_2164; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2233 = wb_state ? _GEN_2212 : _GEN_2176; // @[Conditional.scala 39:67]
  wire  _GEN_2234 = wb_state ? _GEN_2213 : _GEN_2178; // @[Conditional.scala 39:67]
  wire  _GEN_2235 = wb_state ? _GEN_2214 : _GEN_2165; // @[Conditional.scala 39:67]
  wire  _GEN_2236 = wb_state ? _GEN_2215 : _GEN_2179; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2237 = wb_state ? _GEN_2216 : _GEN_2166; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2238 = wb_state ? _GEN_2217 : _GEN_2180; // @[Conditional.scala 39:67]
  wire  _GEN_2239 = wb_state ? _GEN_2218 : _GEN_2182; // @[Conditional.scala 39:67]
  wire  _GEN_2240 = wb_state ? _GEN_2219 : _GEN_2167; // @[Conditional.scala 39:67]
  wire  _GEN_2241 = wb_state ? _GEN_2220 : _GEN_2183; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2242 = wb_state ? _GEN_2221 : _GEN_2168; // @[Conditional.scala 39:67]
  wire [127:0] _GEN_2243 = wb_state ? _GEN_2222 : _GEN_2184; // @[Conditional.scala 39:67]
  wire  _GEN_2244 = wb_state ? _GEN_2223 : _GEN_2186; // @[Conditional.scala 39:67]
  wire  _GEN_2246 = _T_63 ? _GEN_2196 : _GEN_2225; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2247 = _T_63 ? _GEN_2197 : _GEN_2227; // @[Conditional.scala 40:58]
  wire  _GEN_2248 = _T_63 ? _GEN_2198 : _GEN_2230; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2249 = _T_63 ? _GEN_2199 : _GEN_2232; // @[Conditional.scala 40:58]
  wire  _GEN_2250 = _T_63 ? _GEN_2200 : _GEN_2235; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2251 = _T_63 ? _GEN_2201 : _GEN_2237; // @[Conditional.scala 40:58]
  wire  _GEN_2252 = _T_63 ? _GEN_2202 : _GEN_2240; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2253 = _T_63 ? _GEN_2203 : _GEN_2242; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2256 = _T_63 ? _GEN_2162 : _GEN_2227; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2260 = _T_63 ? _GEN_2164 : _GEN_2232; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2264 = _T_63 ? _GEN_2166 : _GEN_2237; // @[Conditional.scala 40:58]
  wire [5:0] _GEN_2268 = _T_63 ? _GEN_2168 : _GEN_2242; // @[Conditional.scala 40:58]
  reg [7:0] counter; // @[Cache_Soc.scala 296:24]
  wire  check_finish = counter == 8'hff; // @[Cache_Soc.scala 297:30]
  wire [5:0] tag_counter = counter[7:2]; // @[Cache_Soc.scala 298:28]
  wire [1:0] way_counter = counter[1:0]; // @[Cache_Soc.scala 299:28]
  wire  _T_73 = 3'h0 == fence_state; // @[Conditional.scala 37:30]
  wire  _T_74 = 3'h1 == fence_state; // @[Conditional.scala 37:30]
  wire  _T_78 = 3'h2 == fence_state; // @[Conditional.scala 37:30]
  wire  _T_79 = way_counter == 2'h0; // @[Cache_Soc.scala 316:27]
  wire [5:0] _GEN_2272 = way_counter == 2'h0 ? tag_counter : _GEN_2256; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 317:28]
  wire [5:0] _GEN_2274 = _T_79 ? tag_counter : _GEN_2247; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2275 = _T_79 | _GEN_2246; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire  _T_81 = way_counter == 2'h1; // @[Cache_Soc.scala 324:31]
  wire [5:0] _GEN_2276 = way_counter == 2'h1 ? tag_counter : _GEN_2249; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2277 = way_counter == 2'h1 | _GEN_2248; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire  _T_82 = way_counter == 2'h2; // @[Cache_Soc.scala 324:31]
  wire [5:0] _GEN_2278 = way_counter == 2'h2 ? tag_counter : _GEN_2251; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2279 = way_counter == 2'h2 | _GEN_2250; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire  _T_83 = way_counter == 2'h3; // @[Cache_Soc.scala 324:31]
  wire [5:0] _GEN_2280 = way_counter == 2'h3 ? tag_counter : _GEN_2253; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2281 = way_counter == 2'h3 | _GEN_2252; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [7:0] _counter_T_1 = counter + 8'h1; // @[Cache_Soc.scala 330:30]
  wire [2:0] _fence_state_T = check_finish ? 3'h5 : 3'h2; // @[Cache_Soc.scala 331:29]
  wire  _GEN_2293 = _T_81 ? meta_1_io_fence_dirty : way_counter == 2'h0 & meta_0_io_fence_dirty; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 318:20]
  wire  _GEN_2313 = _T_82 ? meta_2_io_fence_dirty : _GEN_2293; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 318:20]
  wire  _GEN_2333 = _T_83 ? meta_3_io_fence_dirty : _GEN_2313; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 318:20]
  wire  _GEN_2399 = _T_74 ? 1'h0 : _T_78 & _GEN_2333; // @[Conditional.scala 39:67]
  wire  is_dirty = _T_73 ? 1'h0 : _GEN_2399; // @[Conditional.scala 40:58]
  wire [2:0] _GEN_2282 = is_dirty ? 3'h3 : _fence_state_T; // @[Cache_Soc.scala 321:25 Cache_Soc.scala 322:23 Cache_Soc.scala 331:23]
  wire [5:0] _GEN_2283 = is_dirty ? _GEN_2274 : _GEN_2247; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2284 = is_dirty ? _GEN_2275 : _GEN_2246; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2285 = is_dirty ? _GEN_2276 : _GEN_2249; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2286 = is_dirty ? _GEN_2277 : _GEN_2248; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2287 = is_dirty ? _GEN_2278 : _GEN_2251; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2288 = is_dirty ? _GEN_2279 : _GEN_2250; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2289 = is_dirty ? _GEN_2280 : _GEN_2253; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2290 = is_dirty ? _GEN_2281 : _GEN_2252; // @[Cache_Soc.scala 321:25]
  wire [7:0] _GEN_2291 = is_dirty ? counter : _counter_T_1; // @[Cache_Soc.scala 321:25 Cache_Soc.scala 296:24 Cache_Soc.scala 330:19]
  wire [5:0] _GEN_2292 = _T_81 ? tag_counter : _GEN_2260; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 317:28]
  wire [5:0] _GEN_2294 = _T_79 ? tag_counter : _GEN_2283; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2295 = _T_79 | _GEN_2284; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2296 = way_counter == 2'h1 ? tag_counter : _GEN_2285; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2297 = way_counter == 2'h1 | _GEN_2286; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2298 = way_counter == 2'h2 ? tag_counter : _GEN_2287; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2299 = way_counter == 2'h2 | _GEN_2288; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2300 = way_counter == 2'h3 ? tag_counter : _GEN_2289; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2301 = way_counter == 2'h3 | _GEN_2290; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2303 = is_dirty ? _GEN_2294 : _GEN_2283; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2304 = is_dirty ? _GEN_2295 : _GEN_2284; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2305 = is_dirty ? _GEN_2296 : _GEN_2285; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2306 = is_dirty ? _GEN_2297 : _GEN_2286; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2307 = is_dirty ? _GEN_2298 : _GEN_2287; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2308 = is_dirty ? _GEN_2299 : _GEN_2288; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2309 = is_dirty ? _GEN_2300 : _GEN_2289; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2310 = is_dirty ? _GEN_2301 : _GEN_2290; // @[Cache_Soc.scala 321:25]
  wire [7:0] _GEN_2311 = is_dirty ? _GEN_2291 : _counter_T_1; // @[Cache_Soc.scala 321:25 Cache_Soc.scala 330:19]
  wire [5:0] _GEN_2312 = _T_82 ? tag_counter : _GEN_2264; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 317:28]
  wire [5:0] _GEN_2314 = _T_79 ? tag_counter : _GEN_2303; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2315 = _T_79 | _GEN_2304; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2316 = way_counter == 2'h1 ? tag_counter : _GEN_2305; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2317 = way_counter == 2'h1 | _GEN_2306; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2318 = way_counter == 2'h2 ? tag_counter : _GEN_2307; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2319 = way_counter == 2'h2 | _GEN_2308; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2320 = way_counter == 2'h3 ? tag_counter : _GEN_2309; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2321 = way_counter == 2'h3 | _GEN_2310; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2323 = is_dirty ? _GEN_2314 : _GEN_2303; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2324 = is_dirty ? _GEN_2315 : _GEN_2304; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2325 = is_dirty ? _GEN_2316 : _GEN_2305; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2326 = is_dirty ? _GEN_2317 : _GEN_2306; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2327 = is_dirty ? _GEN_2318 : _GEN_2307; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2328 = is_dirty ? _GEN_2319 : _GEN_2308; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2329 = is_dirty ? _GEN_2320 : _GEN_2309; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2330 = is_dirty ? _GEN_2321 : _GEN_2310; // @[Cache_Soc.scala 321:25]
  wire [7:0] _GEN_2331 = is_dirty ? _GEN_2311 : _counter_T_1; // @[Cache_Soc.scala 321:25 Cache_Soc.scala 330:19]
  wire [5:0] _GEN_2332 = _T_83 ? tag_counter : _GEN_2268; // @[Cache_Soc.scala 316:36 Cache_Soc.scala 317:28]
  wire [5:0] _GEN_2334 = _T_79 ? tag_counter : _GEN_2323; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2335 = _T_79 | _GEN_2324; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2336 = way_counter == 2'h1 ? tag_counter : _GEN_2325; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2337 = way_counter == 2'h1 | _GEN_2326; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2338 = way_counter == 2'h2 ? tag_counter : _GEN_2327; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2339 = way_counter == 2'h2 | _GEN_2328; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2340 = way_counter == 2'h3 ? tag_counter : _GEN_2329; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 325:28]
  wire  _GEN_2341 = way_counter == 2'h3 | _GEN_2330; // @[Cache_Soc.scala 324:40 Cache_Soc.scala 326:26]
  wire [5:0] _GEN_2343 = is_dirty ? _GEN_2334 : _GEN_2323; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2344 = is_dirty ? _GEN_2335 : _GEN_2324; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2345 = is_dirty ? _GEN_2336 : _GEN_2325; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2346 = is_dirty ? _GEN_2337 : _GEN_2326; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2347 = is_dirty ? _GEN_2338 : _GEN_2327; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2348 = is_dirty ? _GEN_2339 : _GEN_2328; // @[Cache_Soc.scala 321:25]
  wire [5:0] _GEN_2349 = is_dirty ? _GEN_2340 : _GEN_2329; // @[Cache_Soc.scala 321:25]
  wire  _GEN_2350 = is_dirty ? _GEN_2341 : _GEN_2330; // @[Cache_Soc.scala 321:25]
  wire [7:0] _GEN_2351 = is_dirty ? _GEN_2331 : _counter_T_1; // @[Cache_Soc.scala 321:25 Cache_Soc.scala 330:19]
  wire  _T_99 = 3'h3 == fence_state; // @[Conditional.scala 37:30]
  wire [21:0] _GEN_2353 = 2'h1 == way_counter ? tag_1 : tag_0; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_2354 = 2'h2 == way_counter ? tag_2 : _GEN_2353; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [21:0] _GEN_2355 = 2'h3 == way_counter ? tag_3 : _GEN_2354; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _io_out_wr_addr_T_3 = {_GEN_2355,tag_counter,4'h0}; // @[Cat.scala 30:58]
  wire [127:0] _GEN_2357 = 2'h1 == way_counter ? io_sram_1_rdata : io_sram_0_rdata; // @[Cache_Soc.scala 340:19 Cache_Soc.scala 340:19]
  wire [127:0] _GEN_2358 = 2'h2 == way_counter ? io_sram_2_rdata : _GEN_2357; // @[Cache_Soc.scala 340:19 Cache_Soc.scala 340:19]
  wire [127:0] _GEN_2359 = 2'h3 == way_counter ? io_sram_3_rdata : _GEN_2358; // @[Cache_Soc.scala 340:19 Cache_Soc.scala 340:19]
  wire [2:0] _GEN_2360 = _T_33 ? 3'h4 : fence_state; // @[Cache_Soc.scala 341:39 Cache_Soc.scala 342:21 Cache_Soc.scala 43:28]
  wire  _T_101 = 3'h4 == fence_state; // @[Conditional.scala 37:30]
  wire [7:0] _GEN_2361 = io_out_wr_ok ? _counter_T_1 : counter; // @[Cache_Soc.scala 346:24 Cache_Soc.scala 347:17 Cache_Soc.scala 296:24]
  wire [2:0] _GEN_2362 = io_out_wr_ok ? _fence_state_T : fence_state; // @[Cache_Soc.scala 346:24 Cache_Soc.scala 348:21 Cache_Soc.scala 43:28]
  wire  _T_102 = 3'h5 == fence_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_2364 = _T_102 ? 3'h0 : fence_state; // @[Conditional.scala 39:67 Cache_Soc.scala 356:19 Cache_Soc.scala 43:28]
  wire [7:0] _GEN_2365 = _T_101 ? _GEN_2361 : counter; // @[Conditional.scala 39:67 Cache_Soc.scala 296:24]
  wire [2:0] _GEN_2366 = _T_101 ? _GEN_2362 : _GEN_2364; // @[Conditional.scala 39:67]
  wire  _GEN_2367 = _T_101 ? 1'h0 : _T_102; // @[Conditional.scala 39:67 Cache_Soc.scala 34:16]
  wire  _GEN_2368 = _T_99 | _GEN_2169; // @[Conditional.scala 39:67 Cache_Soc.scala 336:18]
  wire [2:0] _GEN_2369 = _T_99 ? 3'h3 : _io_out_wr_size_T; // @[Conditional.scala 39:67 Cache_Soc.scala 337:19 Cache_Soc.scala 176:15]
  wire [31:0] _GEN_2370 = _T_99 ? _io_out_wr_addr_T_3 : _io_out_wr_addr_T_2; // @[Conditional.scala 39:67 Cache_Soc.scala 338:19 Cache_Soc.scala 177:15]
  wire [7:0] _GEN_2371 = _T_99 ? 8'hff : _io_out_wr_wstrb_T; // @[Conditional.scala 39:67 Cache_Soc.scala 339:20 Cache_Soc.scala 178:16]
  wire [127:0] _GEN_2372 = _T_99 ? _GEN_2359 : _io_out_wr_data_T_1; // @[Conditional.scala 39:67 Cache_Soc.scala 340:19 Cache_Soc.scala 179:15]
  wire [2:0] _GEN_2373 = _T_99 ? _GEN_2360 : _GEN_2366; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_2374 = _T_99 ? counter : _GEN_2365; // @[Conditional.scala 39:67 Cache_Soc.scala 296:24]
  wire  _GEN_2375 = _T_99 ? 1'h0 : _GEN_2367; // @[Conditional.scala 39:67 Cache_Soc.scala 34:16]
  wire [5:0] _GEN_2376 = _T_78 ? _GEN_2272 : _GEN_2256; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2379 = _T_78 ? _GEN_2343 : _GEN_2247; // @[Conditional.scala 39:67]
  wire  _GEN_2380 = _T_78 ? _GEN_2344 : _GEN_2246; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2381 = _T_78 ? _GEN_2345 : _GEN_2249; // @[Conditional.scala 39:67]
  wire  _GEN_2382 = _T_78 ? _GEN_2346 : _GEN_2248; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2383 = _T_78 ? _GEN_2347 : _GEN_2251; // @[Conditional.scala 39:67]
  wire  _GEN_2384 = _T_78 ? _GEN_2348 : _GEN_2250; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2385 = _T_78 ? _GEN_2349 : _GEN_2253; // @[Conditional.scala 39:67]
  wire  _GEN_2386 = _T_78 ? _GEN_2350 : _GEN_2252; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2388 = _T_78 ? _GEN_2292 : _GEN_2260; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2389 = _T_78 ? _GEN_2312 : _GEN_2264; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2390 = _T_78 ? _GEN_2332 : _GEN_2268; // @[Conditional.scala 39:67]
  wire  _GEN_2391 = _T_78 ? _GEN_2169 : _GEN_2368; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2392 = _T_78 ? _io_out_wr_size_T : _GEN_2369; // @[Conditional.scala 39:67 Cache_Soc.scala 176:15]
  wire [31:0] _GEN_2393 = _T_78 ? _io_out_wr_addr_T_2 : _GEN_2370; // @[Conditional.scala 39:67 Cache_Soc.scala 177:15]
  wire [7:0] _GEN_2394 = _T_78 ? _io_out_wr_wstrb_T : _GEN_2371; // @[Conditional.scala 39:67 Cache_Soc.scala 178:16]
  wire [127:0] _GEN_2395 = _T_78 ? _io_out_wr_data_T_1 : _GEN_2372; // @[Conditional.scala 39:67 Cache_Soc.scala 179:15]
  wire  _GEN_2396 = _T_78 ? 1'h0 : _GEN_2375; // @[Conditional.scala 39:67 Cache_Soc.scala 34:16]
  wire [5:0] _GEN_2398 = _T_74 ? _GEN_2256 : _GEN_2376; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2400 = _T_74 ? _GEN_2247 : _GEN_2379; // @[Conditional.scala 39:67]
  wire  _GEN_2401 = _T_74 ? _GEN_2246 : _GEN_2380; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2402 = _T_74 ? _GEN_2249 : _GEN_2381; // @[Conditional.scala 39:67]
  wire  _GEN_2403 = _T_74 ? _GEN_2248 : _GEN_2382; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2404 = _T_74 ? _GEN_2251 : _GEN_2383; // @[Conditional.scala 39:67]
  wire  _GEN_2405 = _T_74 ? _GEN_2250 : _GEN_2384; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2406 = _T_74 ? _GEN_2253 : _GEN_2385; // @[Conditional.scala 39:67]
  wire  _GEN_2407 = _T_74 ? _GEN_2252 : _GEN_2386; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2409 = _T_74 ? _GEN_2260 : _GEN_2388; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2410 = _T_74 ? _GEN_2264 : _GEN_2389; // @[Conditional.scala 39:67]
  wire [5:0] _GEN_2411 = _T_74 ? _GEN_2268 : _GEN_2390; // @[Conditional.scala 39:67]
  wire  _GEN_2412 = _T_74 ? _GEN_2169 : _GEN_2391; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2413 = _T_74 ? _io_out_wr_size_T : _GEN_2392; // @[Conditional.scala 39:67 Cache_Soc.scala 176:15]
  wire [31:0] _GEN_2414 = _T_74 ? _io_out_wr_addr_T_2 : _GEN_2393; // @[Conditional.scala 39:67 Cache_Soc.scala 177:15]
  wire [7:0] _GEN_2415 = _T_74 ? _io_out_wr_wstrb_T : _GEN_2394; // @[Conditional.scala 39:67 Cache_Soc.scala 178:16]
  wire [127:0] _GEN_2416 = _T_74 ? _io_out_wr_data_T_1 : _GEN_2395; // @[Conditional.scala 39:67 Cache_Soc.scala 179:15]
  wire  _GEN_2417 = _T_74 ? 1'h0 : _GEN_2396; // @[Conditional.scala 39:67 Cache_Soc.scala 34:16]
  META meta_0 ( // @[Cache_Soc.scala 24:22]
    .clock(meta_0_clock),
    .reset(meta_0_reset),
    .io_index(meta_0_io_index),
    .io_tag_r(meta_0_io_tag_r),
    .io_tag_w(meta_0_io_tag_w),
    .io_tag_wen(meta_0_io_tag_wen),
    .io_dirty_r(meta_0_io_dirty_r),
    .io_dirty_w(meta_0_io_dirty_w),
    .io_dirty_wen(meta_0_io_dirty_wen),
    .io_valid_r(meta_0_io_valid_r),
    .io_fence(meta_0_io_fence),
    .io_fence_dirty(meta_0_io_fence_dirty)
  );
  META meta_1 ( // @[Cache_Soc.scala 24:22]
    .clock(meta_1_clock),
    .reset(meta_1_reset),
    .io_index(meta_1_io_index),
    .io_tag_r(meta_1_io_tag_r),
    .io_tag_w(meta_1_io_tag_w),
    .io_tag_wen(meta_1_io_tag_wen),
    .io_dirty_r(meta_1_io_dirty_r),
    .io_dirty_w(meta_1_io_dirty_w),
    .io_dirty_wen(meta_1_io_dirty_wen),
    .io_valid_r(meta_1_io_valid_r),
    .io_fence(meta_1_io_fence),
    .io_fence_dirty(meta_1_io_fence_dirty)
  );
  META meta_2 ( // @[Cache_Soc.scala 24:22]
    .clock(meta_2_clock),
    .reset(meta_2_reset),
    .io_index(meta_2_io_index),
    .io_tag_r(meta_2_io_tag_r),
    .io_tag_w(meta_2_io_tag_w),
    .io_tag_wen(meta_2_io_tag_wen),
    .io_dirty_r(meta_2_io_dirty_r),
    .io_dirty_w(meta_2_io_dirty_w),
    .io_dirty_wen(meta_2_io_dirty_wen),
    .io_valid_r(meta_2_io_valid_r),
    .io_fence(meta_2_io_fence),
    .io_fence_dirty(meta_2_io_fence_dirty)
  );
  META meta_3 ( // @[Cache_Soc.scala 24:22]
    .clock(meta_3_clock),
    .reset(meta_3_reset),
    .io_index(meta_3_io_index),
    .io_tag_r(meta_3_io_tag_r),
    .io_tag_w(meta_3_io_tag_w),
    .io_tag_wen(meta_3_io_tag_wen),
    .io_dirty_r(meta_3_io_dirty_r),
    .io_dirty_w(meta_3_io_dirty_w),
    .io_dirty_wen(meta_3_io_dirty_wen),
    .io_valid_r(meta_3_io_valid_r),
    .io_fence(meta_3_io_fence),
    .io_fence_dirty(meta_3_io_fence_dirty)
  );
  assign io_in_fence_finish = _T_73 ? 1'h0 : _GEN_2417; // @[Conditional.scala 40:58 Cache_Soc.scala 34:16]
  assign io_in_data_ok = _T_1 | _T_2 & (rb_uncache & rb_op & io_out_wr_ok | io_out_ret_valid); // @[Cache_Soc.scala 157:51]
  assign io_in_rdata = _T_1 ? load_res : _io_in_rdata_T_4; // @[Cache_Soc.scala 170:18]
  assign io_in_inst = _T_1 ? load_inst : _io_in_inst_T_4; // @[Cache_Soc.scala 171:17]
  assign io_out_rd_req = _T_18 ? 1'h0 : _GEN_2143; // @[Conditional.scala 40:58 Cache_Soc.scala 174:14]
  assign io_out_rd_size = rb_uncache ? 3'h2 : 3'h3; // @[Cache_Soc.scala 181:21]
  assign io_out_rd_addr = rb_uncache ? _io_out_wr_addr_T : _io_out_rd_addr_T_1; // @[Cache_Soc.scala 182:21]
  assign io_out_wr_req = _T_73 ? _GEN_2169 : _GEN_2412; // @[Conditional.scala 40:58]
  assign io_out_wr_size = _T_73 ? _io_out_wr_size_T : _GEN_2413; // @[Conditional.scala 40:58 Cache_Soc.scala 176:15]
  assign io_out_wr_addr = _T_73 ? _io_out_wr_addr_T_2 : _GEN_2414; // @[Conditional.scala 40:58 Cache_Soc.scala 177:15]
  assign io_out_wr_wstrb = _T_73 ? _io_out_wr_wstrb_T : _GEN_2415; // @[Conditional.scala 40:58 Cache_Soc.scala 178:16]
  assign io_out_wr_data = _T_73 ? _io_out_wr_data_T_1 : _GEN_2416; // @[Conditional.scala 40:58 Cache_Soc.scala 179:15]
  assign io_sram_0_en = _T_73 ? _GEN_2246 : _GEN_2401; // @[Conditional.scala 40:58]
  assign io_sram_0_wen = _T_63 ? _GEN_2171 : _GEN_2226; // @[Conditional.scala 40:58]
  assign io_sram_0_addr = _T_73 ? _GEN_2247 : _GEN_2400; // @[Conditional.scala 40:58]
  assign io_sram_0_wdata = _T_63 ? _GEN_2172 : _GEN_2228; // @[Conditional.scala 40:58]
  assign io_sram_1_en = _T_73 ? _GEN_2248 : _GEN_2403; // @[Conditional.scala 40:58]
  assign io_sram_1_wen = _T_63 ? _GEN_2175 : _GEN_2231; // @[Conditional.scala 40:58]
  assign io_sram_1_addr = _T_73 ? _GEN_2249 : _GEN_2402; // @[Conditional.scala 40:58]
  assign io_sram_1_wdata = _T_63 ? _GEN_2176 : _GEN_2233; // @[Conditional.scala 40:58]
  assign io_sram_2_en = _T_73 ? _GEN_2250 : _GEN_2405; // @[Conditional.scala 40:58]
  assign io_sram_2_wen = _T_63 ? _GEN_2179 : _GEN_2236; // @[Conditional.scala 40:58]
  assign io_sram_2_addr = _T_73 ? _GEN_2251 : _GEN_2404; // @[Conditional.scala 40:58]
  assign io_sram_2_wdata = _T_63 ? _GEN_2180 : _GEN_2238; // @[Conditional.scala 40:58]
  assign io_sram_3_en = _T_73 ? _GEN_2252 : _GEN_2407; // @[Conditional.scala 40:58]
  assign io_sram_3_wen = _T_63 ? _GEN_2183 : _GEN_2241; // @[Conditional.scala 40:58]
  assign io_sram_3_addr = _T_73 ? _GEN_2253 : _GEN_2406; // @[Conditional.scala 40:58]
  assign io_sram_3_wdata = _T_63 ? _GEN_2184 : _GEN_2243; // @[Conditional.scala 40:58]
  assign meta_0_clock = clock;
  assign meta_0_reset = reset;
  assign meta_0_io_index = _T_73 ? _GEN_2256 : _GEN_2398; // @[Conditional.scala 40:58]
  assign meta_0_io_tag_w = _T_18 ? 22'h0 : _GEN_2146; // @[Conditional.scala 40:58 Cache_Soc.scala 30:16]
  assign meta_0_io_tag_wen = _T_18 ? 1'h0 : _GEN_2144; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  assign meta_0_io_dirty_w = _T_63 ? _GEN_2174 : _GEN_2229; // @[Conditional.scala 40:58]
  assign meta_0_io_dirty_wen = _T_63 ? _GEN_2171 : _GEN_2226; // @[Conditional.scala 40:58]
  assign meta_0_io_fence = _T_73 ? 1'h0 : _GEN_2417; // @[Conditional.scala 40:58 Cache_Soc.scala 34:16]
  assign meta_1_clock = clock;
  assign meta_1_reset = reset;
  assign meta_1_io_index = _T_73 ? _GEN_2260 : _GEN_2409; // @[Conditional.scala 40:58]
  assign meta_1_io_tag_w = _T_18 ? 22'h0 : _GEN_2150; // @[Conditional.scala 40:58 Cache_Soc.scala 30:16]
  assign meta_1_io_tag_wen = _T_18 ? 1'h0 : _GEN_2148; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  assign meta_1_io_dirty_w = _T_63 ? _GEN_2178 : _GEN_2234; // @[Conditional.scala 40:58]
  assign meta_1_io_dirty_wen = _T_63 ? _GEN_2175 : _GEN_2231; // @[Conditional.scala 40:58]
  assign meta_1_io_fence = _T_73 ? 1'h0 : _GEN_2417; // @[Conditional.scala 40:58 Cache_Soc.scala 34:16]
  assign meta_2_clock = clock;
  assign meta_2_reset = reset;
  assign meta_2_io_index = _T_73 ? _GEN_2264 : _GEN_2410; // @[Conditional.scala 40:58]
  assign meta_2_io_tag_w = _T_18 ? 22'h0 : _GEN_2154; // @[Conditional.scala 40:58 Cache_Soc.scala 30:16]
  assign meta_2_io_tag_wen = _T_18 ? 1'h0 : _GEN_2152; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  assign meta_2_io_dirty_w = _T_63 ? _GEN_2182 : _GEN_2239; // @[Conditional.scala 40:58]
  assign meta_2_io_dirty_wen = _T_63 ? _GEN_2179 : _GEN_2236; // @[Conditional.scala 40:58]
  assign meta_2_io_fence = _T_73 ? 1'h0 : _GEN_2417; // @[Conditional.scala 40:58 Cache_Soc.scala 34:16]
  assign meta_3_clock = clock;
  assign meta_3_reset = reset;
  assign meta_3_io_index = _T_73 ? _GEN_2268 : _GEN_2411; // @[Conditional.scala 40:58]
  assign meta_3_io_tag_w = _T_18 ? 22'h0 : _GEN_2158; // @[Conditional.scala 40:58 Cache_Soc.scala 30:16]
  assign meta_3_io_tag_wen = _T_18 ? 1'h0 : _GEN_2156; // @[Conditional.scala 40:58 Cache_Soc.scala 18:11]
  assign meta_3_io_dirty_w = _T_63 ? _GEN_2186 : _GEN_2244; // @[Conditional.scala 40:58]
  assign meta_3_io_dirty_wen = _T_63 ? _GEN_2183 : _GEN_2241; // @[Conditional.scala 40:58]
  assign meta_3_io_fence = _T_73 ? 1'h0 : _GEN_2417; // @[Conditional.scala 40:58 Cache_Soc.scala 34:16]
  always @(posedge clock) begin
    if (reset) begin // @[Cache_Soc.scala 41:22]
      state <= 3'h0; // @[Cache_Soc.scala 41:22]
    end else if (_T_18) begin // @[Conditional.scala 40:58]
      if (_T_10) begin // @[Cache_Soc.scala 186:34]
        state <= 3'h1; // @[Cache_Soc.scala 187:15]
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      if (cache_hit & _T_10) begin // @[Cache_Soc.scala 198:49]
        state <= 3'h1; // @[Cache_Soc.scala 199:15]
      end else begin
        state <= _GEN_2032;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      state <= _GEN_2037;
    end else begin
      state <= _GEN_2089;
    end
    if (reset) begin // @[Cache_Soc.scala 42:25]
      wb_state <= 1'h0; // @[Cache_Soc.scala 42:25]
    end else if (_T_63) begin // @[Conditional.scala 40:58]
      wb_state <= _GEN_2195;
    end else if (wb_state) begin // @[Conditional.scala 39:67]
      wb_state <= 1'h0; // @[Cache_Soc.scala 278:16]
    end
    if (reset) begin // @[Cache_Soc.scala 43:28]
      fence_state <= 3'h0; // @[Cache_Soc.scala 43:28]
    end else if (_T_73) begin // @[Conditional.scala 40:58]
      if (io_in_fence) begin // @[Cache_Soc.scala 305:23]
        fence_state <= 3'h1; // @[Cache_Soc.scala 306:21]
      end
    end else if (_T_74) begin // @[Conditional.scala 39:67]
      if (_addr_ok_T & _T_63) begin // @[Cache_Soc.scala 310:57]
        fence_state <= 3'h2; // @[Cache_Soc.scala 311:21]
      end
    end else if (_T_78) begin // @[Conditional.scala 39:67]
      fence_state <= _GEN_2282;
    end else begin
      fence_state <= _GEN_2373;
    end
    if (reset) begin // @[Cache_Soc.scala 55:22]
      rb_op <= 1'h0; // @[Cache_Soc.scala 55:22]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_op <= io_in_op; // @[Cache_Soc.scala 128:11]
    end
    if (reset) begin // @[Cache_Soc.scala 56:27]
      rb_uncache <= 1'h0; // @[Cache_Soc.scala 56:27]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_uncache <= in_uncache; // @[Cache_Soc.scala 129:16]
    end
    if (reset) begin // @[Cache_Soc.scala 57:25]
      rb_index <= 6'h0; // @[Cache_Soc.scala 57:25]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_index <= in_index; // @[Cache_Soc.scala 130:14]
    end
    if (reset) begin // @[Cache_Soc.scala 58:23]
      rb_tag <= 22'h0; // @[Cache_Soc.scala 58:23]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_tag <= in_tag; // @[Cache_Soc.scala 131:12]
    end
    if (reset) begin // @[Cache_Soc.scala 59:26]
      rb_offset <= 4'h0; // @[Cache_Soc.scala 59:26]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_offset <= in_offset; // @[Cache_Soc.scala 132:15]
    end
    if (reset) begin // @[Cache_Soc.scala 60:25]
      rb_wstrb <= 8'h0; // @[Cache_Soc.scala 60:25]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_wstrb <= io_in_wstrb; // @[Cache_Soc.scala 133:14]
    end
    if (reset) begin // @[Cache_Soc.scala 61:25]
      rb_wdata <= 64'h0; // @[Cache_Soc.scala 61:25]
    end else if (io_in_valid & addr_ok) begin // @[Cache_Soc.scala 127:30]
      rb_wdata <= io_in_wdata; // @[Cache_Soc.scala 134:14]
    end
    if (reset) begin // @[Cache_Soc.scala 64:26]
      wb_hitway <= 2'h0; // @[Cache_Soc.scala 64:26]
    end else if (_T_1 & rb_op) begin // @[Cache_Soc.scala 138:61]
      wb_hitway <= _wb_hitway_T_2; // @[Cache_Soc.scala 139:15]
    end
    if (reset) begin // @[Cache_Soc.scala 65:25]
      wb_index <= 6'h0; // @[Cache_Soc.scala 65:25]
    end else if (_T_1 & rb_op) begin // @[Cache_Soc.scala 138:61]
      wb_index <= rb_index; // @[Cache_Soc.scala 140:14]
    end
    if (reset) begin // @[Cache_Soc.scala 67:26]
      wb_offset <= 4'h0; // @[Cache_Soc.scala 67:26]
    end else if (_T_1 & rb_op) begin // @[Cache_Soc.scala 138:61]
      wb_offset <= rb_offset; // @[Cache_Soc.scala 142:15]
    end
    if (reset) begin // @[Cache_Soc.scala 68:25]
      wb_wstrb <= 8'h0; // @[Cache_Soc.scala 68:25]
    end else if (_T_1 & rb_op) begin // @[Cache_Soc.scala 138:61]
      wb_wstrb <= rb_wstrb; // @[Cache_Soc.scala 143:14]
    end
    if (reset) begin // @[Cache_Soc.scala 69:25]
      wb_wdata <= 64'h0; // @[Cache_Soc.scala 69:25]
    end else if (_T_1 & rb_op) begin // @[Cache_Soc.scala 138:61]
      wb_wdata <= rb_wdata; // @[Cache_Soc.scala 144:14]
    end
    if (reset) begin // @[Cache_Soc.scala 72:30]
      replace_valid <= 1'h0; // @[Cache_Soc.scala 72:30]
    end else if (_T & ~cache_hit) begin // @[Cache_Soc.scala 148:41]
      if (2'h3 == replace_way) begin // @[Cache_Soc.scala 149:19]
        replace_valid <= valid_3; // @[Cache_Soc.scala 149:19]
      end else if (2'h2 == replace_way) begin // @[Cache_Soc.scala 149:19]
        replace_valid <= valid_2; // @[Cache_Soc.scala 149:19]
      end else begin
        replace_valid <= _GEN_1998;
      end
    end
    if (reset) begin // @[Cache_Soc.scala 73:30]
      replace_dirty <= 1'h0; // @[Cache_Soc.scala 73:30]
    end else if (_T & ~cache_hit) begin // @[Cache_Soc.scala 148:41]
      if (2'h3 == replace_way) begin // @[Cache_Soc.scala 150:19]
        replace_dirty <= dirty_3; // @[Cache_Soc.scala 150:19]
      end else if (2'h2 == replace_way) begin // @[Cache_Soc.scala 150:19]
        replace_dirty <= dirty_2; // @[Cache_Soc.scala 150:19]
      end else begin
        replace_dirty <= _GEN_2002;
      end
    end
    if (reset) begin // @[Cache_Soc.scala 74:28]
      replace_tag <= 22'h0; // @[Cache_Soc.scala 74:28]
    end else if (_T & ~cache_hit) begin // @[Cache_Soc.scala 148:41]
      if (2'h3 == replace_way) begin // @[Cache_Soc.scala 151:17]
        replace_tag <= tag_3; // @[Cache_Soc.scala 151:17]
      end else if (2'h2 == replace_way) begin // @[Cache_Soc.scala 151:17]
        replace_tag <= tag_2; // @[Cache_Soc.scala 151:17]
      end else begin
        replace_tag <= _GEN_2006;
      end
    end
    if (reset) begin // @[Cache_Soc.scala 75:29]
      replace_data <= 128'h0; // @[Cache_Soc.scala 75:29]
    end else if (_T & ~cache_hit) begin // @[Cache_Soc.scala 148:41]
      if (2'h3 == replace_way) begin // @[Cache_Soc.scala 152:18]
        replace_data <= io_sram_3_rdata; // @[Cache_Soc.scala 152:18]
      end else if (2'h2 == replace_way) begin // @[Cache_Soc.scala 152:18]
        replace_data <= io_sram_2_rdata; // @[Cache_Soc.scala 152:18]
      end else begin
        replace_data <= _GEN_2010;
      end
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_0 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h0 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_0 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_0 <= _GEN_704;
      end
    end else begin
      plru0_0 <= _GEN_704;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_1 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_1 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_1 <= _GEN_705;
      end
    end else begin
      plru0_1 <= _GEN_705;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_2 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_2 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_2 <= _GEN_706;
      end
    end else begin
      plru0_2 <= _GEN_706;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_3 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_3 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_3 <= _GEN_707;
      end
    end else begin
      plru0_3 <= _GEN_707;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_4 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h4 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_4 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_4 <= _GEN_708;
      end
    end else begin
      plru0_4 <= _GEN_708;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_5 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h5 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_5 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_5 <= _GEN_709;
      end
    end else begin
      plru0_5 <= _GEN_709;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_6 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h6 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_6 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_6 <= _GEN_710;
      end
    end else begin
      plru0_6 <= _GEN_710;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_7 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h7 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_7 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_7 <= _GEN_711;
      end
    end else begin
      plru0_7 <= _GEN_711;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_8 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h8 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_8 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_8 <= _GEN_712;
      end
    end else begin
      plru0_8 <= _GEN_712;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_9 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h9 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_9 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_9 <= _GEN_713;
      end
    end else begin
      plru0_9 <= _GEN_713;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_10 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'ha == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_10 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_10 <= _GEN_714;
      end
    end else begin
      plru0_10 <= _GEN_714;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_11 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'hb == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_11 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_11 <= _GEN_715;
      end
    end else begin
      plru0_11 <= _GEN_715;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_12 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'hc == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_12 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_12 <= _GEN_716;
      end
    end else begin
      plru0_12 <= _GEN_716;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_13 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'hd == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_13 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_13 <= _GEN_717;
      end
    end else begin
      plru0_13 <= _GEN_717;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_14 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'he == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_14 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_14 <= _GEN_718;
      end
    end else begin
      plru0_14 <= _GEN_718;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_15 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'hf == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_15 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_15 <= _GEN_719;
      end
    end else begin
      plru0_15 <= _GEN_719;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_16 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h10 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_16 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_16 <= _GEN_720;
      end
    end else begin
      plru0_16 <= _GEN_720;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_17 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h11 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_17 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_17 <= _GEN_721;
      end
    end else begin
      plru0_17 <= _GEN_721;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_18 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h12 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_18 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_18 <= _GEN_722;
      end
    end else begin
      plru0_18 <= _GEN_722;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_19 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h13 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_19 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_19 <= _GEN_723;
      end
    end else begin
      plru0_19 <= _GEN_723;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_20 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h14 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_20 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_20 <= _GEN_724;
      end
    end else begin
      plru0_20 <= _GEN_724;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_21 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h15 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_21 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_21 <= _GEN_725;
      end
    end else begin
      plru0_21 <= _GEN_725;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_22 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h16 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_22 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_22 <= _GEN_726;
      end
    end else begin
      plru0_22 <= _GEN_726;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_23 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h17 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_23 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_23 <= _GEN_727;
      end
    end else begin
      plru0_23 <= _GEN_727;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_24 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h18 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_24 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_24 <= _GEN_728;
      end
    end else begin
      plru0_24 <= _GEN_728;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_25 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h19 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_25 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_25 <= _GEN_729;
      end
    end else begin
      plru0_25 <= _GEN_729;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_26 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1a == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_26 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_26 <= _GEN_730;
      end
    end else begin
      plru0_26 <= _GEN_730;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_27 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1b == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_27 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_27 <= _GEN_731;
      end
    end else begin
      plru0_27 <= _GEN_731;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_28 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1c == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_28 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_28 <= _GEN_732;
      end
    end else begin
      plru0_28 <= _GEN_732;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_29 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1d == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_29 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_29 <= _GEN_733;
      end
    end else begin
      plru0_29 <= _GEN_733;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_30 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1e == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_30 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_30 <= _GEN_734;
      end
    end else begin
      plru0_30 <= _GEN_734;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_31 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h1f == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_31 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_31 <= _GEN_735;
      end
    end else begin
      plru0_31 <= _GEN_735;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_32 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h20 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_32 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_32 <= _GEN_736;
      end
    end else begin
      plru0_32 <= _GEN_736;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_33 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h21 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_33 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_33 <= _GEN_737;
      end
    end else begin
      plru0_33 <= _GEN_737;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_34 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h22 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_34 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_34 <= _GEN_738;
      end
    end else begin
      plru0_34 <= _GEN_738;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_35 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h23 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_35 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_35 <= _GEN_739;
      end
    end else begin
      plru0_35 <= _GEN_739;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_36 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h24 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_36 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_36 <= _GEN_740;
      end
    end else begin
      plru0_36 <= _GEN_740;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_37 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h25 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_37 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_37 <= _GEN_741;
      end
    end else begin
      plru0_37 <= _GEN_741;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_38 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h26 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_38 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_38 <= _GEN_742;
      end
    end else begin
      plru0_38 <= _GEN_742;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_39 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h27 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_39 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_39 <= _GEN_743;
      end
    end else begin
      plru0_39 <= _GEN_743;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_40 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h28 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_40 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_40 <= _GEN_744;
      end
    end else begin
      plru0_40 <= _GEN_744;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_41 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h29 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_41 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_41 <= _GEN_745;
      end
    end else begin
      plru0_41 <= _GEN_745;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_42 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2a == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_42 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_42 <= _GEN_746;
      end
    end else begin
      plru0_42 <= _GEN_746;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_43 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2b == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_43 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_43 <= _GEN_747;
      end
    end else begin
      plru0_43 <= _GEN_747;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_44 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2c == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_44 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_44 <= _GEN_748;
      end
    end else begin
      plru0_44 <= _GEN_748;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_45 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2d == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_45 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_45 <= _GEN_749;
      end
    end else begin
      plru0_45 <= _GEN_749;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_46 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2e == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_46 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_46 <= _GEN_750;
      end
    end else begin
      plru0_46 <= _GEN_750;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_47 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h2f == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_47 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_47 <= _GEN_751;
      end
    end else begin
      plru0_47 <= _GEN_751;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_48 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h30 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_48 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_48 <= _GEN_752;
      end
    end else begin
      plru0_48 <= _GEN_752;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_49 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h31 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_49 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_49 <= _GEN_753;
      end
    end else begin
      plru0_49 <= _GEN_753;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_50 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h32 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_50 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_50 <= _GEN_754;
      end
    end else begin
      plru0_50 <= _GEN_754;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_51 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h33 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_51 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_51 <= _GEN_755;
      end
    end else begin
      plru0_51 <= _GEN_755;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_52 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h34 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_52 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_52 <= _GEN_756;
      end
    end else begin
      plru0_52 <= _GEN_756;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_53 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h35 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_53 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_53 <= _GEN_757;
      end
    end else begin
      plru0_53 <= _GEN_757;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_54 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h36 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_54 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_54 <= _GEN_758;
      end
    end else begin
      plru0_54 <= _GEN_758;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_55 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h37 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_55 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_55 <= _GEN_759;
      end
    end else begin
      plru0_55 <= _GEN_759;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_56 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h38 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_56 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_56 <= _GEN_760;
      end
    end else begin
      plru0_56 <= _GEN_760;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_57 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h39 == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_57 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_57 <= _GEN_761;
      end
    end else begin
      plru0_57 <= _GEN_761;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_58 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3a == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_58 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_58 <= _GEN_762;
      end
    end else begin
      plru0_58 <= _GEN_762;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_59 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3b == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_59 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_59 <= _GEN_763;
      end
    end else begin
      plru0_59 <= _GEN_763;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_60 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3c == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_60 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_60 <= _GEN_764;
      end
    end else begin
      plru0_60 <= _GEN_764;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_61 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3d == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_61 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_61 <= _GEN_765;
      end
    end else begin
      plru0_61 <= _GEN_765;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_62 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3e == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_62 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_62 <= _GEN_766;
      end
    end else begin
      plru0_62 <= _GEN_766;
    end
    if (reset) begin // @[Cache_Soc.scala 89:22]
      plru0_63 <= 1'h0; // @[Cache_Soc.scala 89:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (6'h3f == rb_index) begin // @[Cache_Soc.scala 107:21]
        plru0_63 <= replace_way == 2'h0 | replace_way == 2'h1; // @[Cache_Soc.scala 107:21]
      end else begin
        plru0_63 <= _GEN_767;
      end
    end else begin
      plru0_63 <= _GEN_767;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_0 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_0 <= _GEN_960;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_0 <= _GEN_1024;
      end else begin
        plru1_0 <= _GEN_768;
      end
    end else begin
      plru1_0 <= _GEN_768;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_1 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_1 <= _GEN_961;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_1 <= _GEN_1025;
      end else begin
        plru1_1 <= _GEN_769;
      end
    end else begin
      plru1_1 <= _GEN_769;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_2 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_2 <= _GEN_962;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_2 <= _GEN_1026;
      end else begin
        plru1_2 <= _GEN_770;
      end
    end else begin
      plru1_2 <= _GEN_770;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_3 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_3 <= _GEN_963;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_3 <= _GEN_1027;
      end else begin
        plru1_3 <= _GEN_771;
      end
    end else begin
      plru1_3 <= _GEN_771;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_4 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_4 <= _GEN_964;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_4 <= _GEN_1028;
      end else begin
        plru1_4 <= _GEN_772;
      end
    end else begin
      plru1_4 <= _GEN_772;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_5 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_5 <= _GEN_965;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_5 <= _GEN_1029;
      end else begin
        plru1_5 <= _GEN_773;
      end
    end else begin
      plru1_5 <= _GEN_773;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_6 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_6 <= _GEN_966;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_6 <= _GEN_1030;
      end else begin
        plru1_6 <= _GEN_774;
      end
    end else begin
      plru1_6 <= _GEN_774;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_7 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_7 <= _GEN_967;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_7 <= _GEN_1031;
      end else begin
        plru1_7 <= _GEN_775;
      end
    end else begin
      plru1_7 <= _GEN_775;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_8 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_8 <= _GEN_968;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_8 <= _GEN_1032;
      end else begin
        plru1_8 <= _GEN_776;
      end
    end else begin
      plru1_8 <= _GEN_776;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_9 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_9 <= _GEN_969;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_9 <= _GEN_1033;
      end else begin
        plru1_9 <= _GEN_777;
      end
    end else begin
      plru1_9 <= _GEN_777;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_10 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_10 <= _GEN_970;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_10 <= _GEN_1034;
      end else begin
        plru1_10 <= _GEN_778;
      end
    end else begin
      plru1_10 <= _GEN_778;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_11 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_11 <= _GEN_971;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_11 <= _GEN_1035;
      end else begin
        plru1_11 <= _GEN_779;
      end
    end else begin
      plru1_11 <= _GEN_779;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_12 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_12 <= _GEN_972;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_12 <= _GEN_1036;
      end else begin
        plru1_12 <= _GEN_780;
      end
    end else begin
      plru1_12 <= _GEN_780;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_13 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_13 <= _GEN_973;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_13 <= _GEN_1037;
      end else begin
        plru1_13 <= _GEN_781;
      end
    end else begin
      plru1_13 <= _GEN_781;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_14 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_14 <= _GEN_974;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_14 <= _GEN_1038;
      end else begin
        plru1_14 <= _GEN_782;
      end
    end else begin
      plru1_14 <= _GEN_782;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_15 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_15 <= _GEN_975;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_15 <= _GEN_1039;
      end else begin
        plru1_15 <= _GEN_783;
      end
    end else begin
      plru1_15 <= _GEN_783;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_16 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_16 <= _GEN_976;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_16 <= _GEN_1040;
      end else begin
        plru1_16 <= _GEN_784;
      end
    end else begin
      plru1_16 <= _GEN_784;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_17 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_17 <= _GEN_977;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_17 <= _GEN_1041;
      end else begin
        plru1_17 <= _GEN_785;
      end
    end else begin
      plru1_17 <= _GEN_785;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_18 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_18 <= _GEN_978;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_18 <= _GEN_1042;
      end else begin
        plru1_18 <= _GEN_786;
      end
    end else begin
      plru1_18 <= _GEN_786;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_19 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_19 <= _GEN_979;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_19 <= _GEN_1043;
      end else begin
        plru1_19 <= _GEN_787;
      end
    end else begin
      plru1_19 <= _GEN_787;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_20 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_20 <= _GEN_980;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_20 <= _GEN_1044;
      end else begin
        plru1_20 <= _GEN_788;
      end
    end else begin
      plru1_20 <= _GEN_788;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_21 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_21 <= _GEN_981;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_21 <= _GEN_1045;
      end else begin
        plru1_21 <= _GEN_789;
      end
    end else begin
      plru1_21 <= _GEN_789;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_22 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_22 <= _GEN_982;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_22 <= _GEN_1046;
      end else begin
        plru1_22 <= _GEN_790;
      end
    end else begin
      plru1_22 <= _GEN_790;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_23 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_23 <= _GEN_983;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_23 <= _GEN_1047;
      end else begin
        plru1_23 <= _GEN_791;
      end
    end else begin
      plru1_23 <= _GEN_791;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_24 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_24 <= _GEN_984;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_24 <= _GEN_1048;
      end else begin
        plru1_24 <= _GEN_792;
      end
    end else begin
      plru1_24 <= _GEN_792;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_25 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_25 <= _GEN_985;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_25 <= _GEN_1049;
      end else begin
        plru1_25 <= _GEN_793;
      end
    end else begin
      plru1_25 <= _GEN_793;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_26 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_26 <= _GEN_986;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_26 <= _GEN_1050;
      end else begin
        plru1_26 <= _GEN_794;
      end
    end else begin
      plru1_26 <= _GEN_794;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_27 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_27 <= _GEN_987;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_27 <= _GEN_1051;
      end else begin
        plru1_27 <= _GEN_795;
      end
    end else begin
      plru1_27 <= _GEN_795;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_28 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_28 <= _GEN_988;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_28 <= _GEN_1052;
      end else begin
        plru1_28 <= _GEN_796;
      end
    end else begin
      plru1_28 <= _GEN_796;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_29 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_29 <= _GEN_989;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_29 <= _GEN_1053;
      end else begin
        plru1_29 <= _GEN_797;
      end
    end else begin
      plru1_29 <= _GEN_797;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_30 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_30 <= _GEN_990;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_30 <= _GEN_1054;
      end else begin
        plru1_30 <= _GEN_798;
      end
    end else begin
      plru1_30 <= _GEN_798;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_31 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_31 <= _GEN_991;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_31 <= _GEN_1055;
      end else begin
        plru1_31 <= _GEN_799;
      end
    end else begin
      plru1_31 <= _GEN_799;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_32 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_32 <= _GEN_992;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_32 <= _GEN_1056;
      end else begin
        plru1_32 <= _GEN_800;
      end
    end else begin
      plru1_32 <= _GEN_800;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_33 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_33 <= _GEN_993;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_33 <= _GEN_1057;
      end else begin
        plru1_33 <= _GEN_801;
      end
    end else begin
      plru1_33 <= _GEN_801;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_34 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_34 <= _GEN_994;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_34 <= _GEN_1058;
      end else begin
        plru1_34 <= _GEN_802;
      end
    end else begin
      plru1_34 <= _GEN_802;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_35 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_35 <= _GEN_995;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_35 <= _GEN_1059;
      end else begin
        plru1_35 <= _GEN_803;
      end
    end else begin
      plru1_35 <= _GEN_803;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_36 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_36 <= _GEN_996;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_36 <= _GEN_1060;
      end else begin
        plru1_36 <= _GEN_804;
      end
    end else begin
      plru1_36 <= _GEN_804;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_37 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_37 <= _GEN_997;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_37 <= _GEN_1061;
      end else begin
        plru1_37 <= _GEN_805;
      end
    end else begin
      plru1_37 <= _GEN_805;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_38 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_38 <= _GEN_998;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_38 <= _GEN_1062;
      end else begin
        plru1_38 <= _GEN_806;
      end
    end else begin
      plru1_38 <= _GEN_806;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_39 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_39 <= _GEN_999;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_39 <= _GEN_1063;
      end else begin
        plru1_39 <= _GEN_807;
      end
    end else begin
      plru1_39 <= _GEN_807;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_40 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_40 <= _GEN_1000;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_40 <= _GEN_1064;
      end else begin
        plru1_40 <= _GEN_808;
      end
    end else begin
      plru1_40 <= _GEN_808;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_41 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_41 <= _GEN_1001;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_41 <= _GEN_1065;
      end else begin
        plru1_41 <= _GEN_809;
      end
    end else begin
      plru1_41 <= _GEN_809;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_42 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_42 <= _GEN_1002;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_42 <= _GEN_1066;
      end else begin
        plru1_42 <= _GEN_810;
      end
    end else begin
      plru1_42 <= _GEN_810;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_43 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_43 <= _GEN_1003;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_43 <= _GEN_1067;
      end else begin
        plru1_43 <= _GEN_811;
      end
    end else begin
      plru1_43 <= _GEN_811;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_44 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_44 <= _GEN_1004;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_44 <= _GEN_1068;
      end else begin
        plru1_44 <= _GEN_812;
      end
    end else begin
      plru1_44 <= _GEN_812;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_45 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_45 <= _GEN_1005;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_45 <= _GEN_1069;
      end else begin
        plru1_45 <= _GEN_813;
      end
    end else begin
      plru1_45 <= _GEN_813;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_46 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_46 <= _GEN_1006;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_46 <= _GEN_1070;
      end else begin
        plru1_46 <= _GEN_814;
      end
    end else begin
      plru1_46 <= _GEN_814;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_47 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_47 <= _GEN_1007;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_47 <= _GEN_1071;
      end else begin
        plru1_47 <= _GEN_815;
      end
    end else begin
      plru1_47 <= _GEN_815;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_48 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_48 <= _GEN_1008;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_48 <= _GEN_1072;
      end else begin
        plru1_48 <= _GEN_816;
      end
    end else begin
      plru1_48 <= _GEN_816;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_49 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_49 <= _GEN_1009;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_49 <= _GEN_1073;
      end else begin
        plru1_49 <= _GEN_817;
      end
    end else begin
      plru1_49 <= _GEN_817;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_50 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_50 <= _GEN_1010;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_50 <= _GEN_1074;
      end else begin
        plru1_50 <= _GEN_818;
      end
    end else begin
      plru1_50 <= _GEN_818;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_51 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_51 <= _GEN_1011;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_51 <= _GEN_1075;
      end else begin
        plru1_51 <= _GEN_819;
      end
    end else begin
      plru1_51 <= _GEN_819;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_52 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_52 <= _GEN_1012;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_52 <= _GEN_1076;
      end else begin
        plru1_52 <= _GEN_820;
      end
    end else begin
      plru1_52 <= _GEN_820;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_53 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_53 <= _GEN_1013;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_53 <= _GEN_1077;
      end else begin
        plru1_53 <= _GEN_821;
      end
    end else begin
      plru1_53 <= _GEN_821;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_54 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_54 <= _GEN_1014;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_54 <= _GEN_1078;
      end else begin
        plru1_54 <= _GEN_822;
      end
    end else begin
      plru1_54 <= _GEN_822;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_55 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_55 <= _GEN_1015;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_55 <= _GEN_1079;
      end else begin
        plru1_55 <= _GEN_823;
      end
    end else begin
      plru1_55 <= _GEN_823;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_56 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_56 <= _GEN_1016;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_56 <= _GEN_1080;
      end else begin
        plru1_56 <= _GEN_824;
      end
    end else begin
      plru1_56 <= _GEN_824;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_57 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_57 <= _GEN_1017;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_57 <= _GEN_1081;
      end else begin
        plru1_57 <= _GEN_825;
      end
    end else begin
      plru1_57 <= _GEN_825;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_58 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_58 <= _GEN_1018;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_58 <= _GEN_1082;
      end else begin
        plru1_58 <= _GEN_826;
      end
    end else begin
      plru1_58 <= _GEN_826;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_59 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_59 <= _GEN_1019;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_59 <= _GEN_1083;
      end else begin
        plru1_59 <= _GEN_827;
      end
    end else begin
      plru1_59 <= _GEN_827;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_60 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_60 <= _GEN_1020;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_60 <= _GEN_1084;
      end else begin
        plru1_60 <= _GEN_828;
      end
    end else begin
      plru1_60 <= _GEN_828;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_61 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_61 <= _GEN_1021;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_61 <= _GEN_1085;
      end else begin
        plru1_61 <= _GEN_829;
      end
    end else begin
      plru1_61 <= _GEN_829;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_62 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_62 <= _GEN_1022;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_62 <= _GEN_1086;
      end else begin
        plru1_62 <= _GEN_830;
      end
    end else begin
      plru1_62 <= _GEN_830;
    end
    if (reset) begin // @[Cache_Soc.scala 90:22]
      plru1_63 <= 1'h0; // @[Cache_Soc.scala 90:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru1_63 <= _GEN_1023;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru1_63 <= _GEN_1087;
      end else begin
        plru1_63 <= _GEN_831;
      end
    end else begin
      plru1_63 <= _GEN_831;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_0 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_0 <= _GEN_832;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_0 <= _GEN_832;
      end else begin
        plru2_0 <= _GEN_1280;
      end
    end else begin
      plru2_0 <= _GEN_832;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_1 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_1 <= _GEN_833;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_1 <= _GEN_833;
      end else begin
        plru2_1 <= _GEN_1281;
      end
    end else begin
      plru2_1 <= _GEN_833;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_2 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_2 <= _GEN_834;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_2 <= _GEN_834;
      end else begin
        plru2_2 <= _GEN_1282;
      end
    end else begin
      plru2_2 <= _GEN_834;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_3 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_3 <= _GEN_835;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_3 <= _GEN_835;
      end else begin
        plru2_3 <= _GEN_1283;
      end
    end else begin
      plru2_3 <= _GEN_835;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_4 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_4 <= _GEN_836;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_4 <= _GEN_836;
      end else begin
        plru2_4 <= _GEN_1284;
      end
    end else begin
      plru2_4 <= _GEN_836;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_5 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_5 <= _GEN_837;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_5 <= _GEN_837;
      end else begin
        plru2_5 <= _GEN_1285;
      end
    end else begin
      plru2_5 <= _GEN_837;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_6 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_6 <= _GEN_838;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_6 <= _GEN_838;
      end else begin
        plru2_6 <= _GEN_1286;
      end
    end else begin
      plru2_6 <= _GEN_838;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_7 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_7 <= _GEN_839;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_7 <= _GEN_839;
      end else begin
        plru2_7 <= _GEN_1287;
      end
    end else begin
      plru2_7 <= _GEN_839;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_8 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_8 <= _GEN_840;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_8 <= _GEN_840;
      end else begin
        plru2_8 <= _GEN_1288;
      end
    end else begin
      plru2_8 <= _GEN_840;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_9 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_9 <= _GEN_841;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_9 <= _GEN_841;
      end else begin
        plru2_9 <= _GEN_1289;
      end
    end else begin
      plru2_9 <= _GEN_841;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_10 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_10 <= _GEN_842;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_10 <= _GEN_842;
      end else begin
        plru2_10 <= _GEN_1290;
      end
    end else begin
      plru2_10 <= _GEN_842;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_11 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_11 <= _GEN_843;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_11 <= _GEN_843;
      end else begin
        plru2_11 <= _GEN_1291;
      end
    end else begin
      plru2_11 <= _GEN_843;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_12 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_12 <= _GEN_844;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_12 <= _GEN_844;
      end else begin
        plru2_12 <= _GEN_1292;
      end
    end else begin
      plru2_12 <= _GEN_844;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_13 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_13 <= _GEN_845;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_13 <= _GEN_845;
      end else begin
        plru2_13 <= _GEN_1293;
      end
    end else begin
      plru2_13 <= _GEN_845;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_14 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_14 <= _GEN_846;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_14 <= _GEN_846;
      end else begin
        plru2_14 <= _GEN_1294;
      end
    end else begin
      plru2_14 <= _GEN_846;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_15 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_15 <= _GEN_847;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_15 <= _GEN_847;
      end else begin
        plru2_15 <= _GEN_1295;
      end
    end else begin
      plru2_15 <= _GEN_847;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_16 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_16 <= _GEN_848;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_16 <= _GEN_848;
      end else begin
        plru2_16 <= _GEN_1296;
      end
    end else begin
      plru2_16 <= _GEN_848;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_17 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_17 <= _GEN_849;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_17 <= _GEN_849;
      end else begin
        plru2_17 <= _GEN_1297;
      end
    end else begin
      plru2_17 <= _GEN_849;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_18 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_18 <= _GEN_850;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_18 <= _GEN_850;
      end else begin
        plru2_18 <= _GEN_1298;
      end
    end else begin
      plru2_18 <= _GEN_850;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_19 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_19 <= _GEN_851;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_19 <= _GEN_851;
      end else begin
        plru2_19 <= _GEN_1299;
      end
    end else begin
      plru2_19 <= _GEN_851;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_20 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_20 <= _GEN_852;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_20 <= _GEN_852;
      end else begin
        plru2_20 <= _GEN_1300;
      end
    end else begin
      plru2_20 <= _GEN_852;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_21 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_21 <= _GEN_853;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_21 <= _GEN_853;
      end else begin
        plru2_21 <= _GEN_1301;
      end
    end else begin
      plru2_21 <= _GEN_853;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_22 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_22 <= _GEN_854;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_22 <= _GEN_854;
      end else begin
        plru2_22 <= _GEN_1302;
      end
    end else begin
      plru2_22 <= _GEN_854;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_23 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_23 <= _GEN_855;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_23 <= _GEN_855;
      end else begin
        plru2_23 <= _GEN_1303;
      end
    end else begin
      plru2_23 <= _GEN_855;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_24 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_24 <= _GEN_856;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_24 <= _GEN_856;
      end else begin
        plru2_24 <= _GEN_1304;
      end
    end else begin
      plru2_24 <= _GEN_856;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_25 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_25 <= _GEN_857;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_25 <= _GEN_857;
      end else begin
        plru2_25 <= _GEN_1305;
      end
    end else begin
      plru2_25 <= _GEN_857;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_26 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_26 <= _GEN_858;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_26 <= _GEN_858;
      end else begin
        plru2_26 <= _GEN_1306;
      end
    end else begin
      plru2_26 <= _GEN_858;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_27 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_27 <= _GEN_859;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_27 <= _GEN_859;
      end else begin
        plru2_27 <= _GEN_1307;
      end
    end else begin
      plru2_27 <= _GEN_859;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_28 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_28 <= _GEN_860;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_28 <= _GEN_860;
      end else begin
        plru2_28 <= _GEN_1308;
      end
    end else begin
      plru2_28 <= _GEN_860;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_29 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_29 <= _GEN_861;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_29 <= _GEN_861;
      end else begin
        plru2_29 <= _GEN_1309;
      end
    end else begin
      plru2_29 <= _GEN_861;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_30 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_30 <= _GEN_862;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_30 <= _GEN_862;
      end else begin
        plru2_30 <= _GEN_1310;
      end
    end else begin
      plru2_30 <= _GEN_862;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_31 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_31 <= _GEN_863;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_31 <= _GEN_863;
      end else begin
        plru2_31 <= _GEN_1311;
      end
    end else begin
      plru2_31 <= _GEN_863;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_32 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_32 <= _GEN_864;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_32 <= _GEN_864;
      end else begin
        plru2_32 <= _GEN_1312;
      end
    end else begin
      plru2_32 <= _GEN_864;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_33 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_33 <= _GEN_865;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_33 <= _GEN_865;
      end else begin
        plru2_33 <= _GEN_1313;
      end
    end else begin
      plru2_33 <= _GEN_865;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_34 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_34 <= _GEN_866;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_34 <= _GEN_866;
      end else begin
        plru2_34 <= _GEN_1314;
      end
    end else begin
      plru2_34 <= _GEN_866;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_35 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_35 <= _GEN_867;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_35 <= _GEN_867;
      end else begin
        plru2_35 <= _GEN_1315;
      end
    end else begin
      plru2_35 <= _GEN_867;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_36 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_36 <= _GEN_868;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_36 <= _GEN_868;
      end else begin
        plru2_36 <= _GEN_1316;
      end
    end else begin
      plru2_36 <= _GEN_868;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_37 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_37 <= _GEN_869;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_37 <= _GEN_869;
      end else begin
        plru2_37 <= _GEN_1317;
      end
    end else begin
      plru2_37 <= _GEN_869;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_38 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_38 <= _GEN_870;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_38 <= _GEN_870;
      end else begin
        plru2_38 <= _GEN_1318;
      end
    end else begin
      plru2_38 <= _GEN_870;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_39 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_39 <= _GEN_871;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_39 <= _GEN_871;
      end else begin
        plru2_39 <= _GEN_1319;
      end
    end else begin
      plru2_39 <= _GEN_871;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_40 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_40 <= _GEN_872;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_40 <= _GEN_872;
      end else begin
        plru2_40 <= _GEN_1320;
      end
    end else begin
      plru2_40 <= _GEN_872;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_41 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_41 <= _GEN_873;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_41 <= _GEN_873;
      end else begin
        plru2_41 <= _GEN_1321;
      end
    end else begin
      plru2_41 <= _GEN_873;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_42 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_42 <= _GEN_874;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_42 <= _GEN_874;
      end else begin
        plru2_42 <= _GEN_1322;
      end
    end else begin
      plru2_42 <= _GEN_874;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_43 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_43 <= _GEN_875;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_43 <= _GEN_875;
      end else begin
        plru2_43 <= _GEN_1323;
      end
    end else begin
      plru2_43 <= _GEN_875;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_44 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_44 <= _GEN_876;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_44 <= _GEN_876;
      end else begin
        plru2_44 <= _GEN_1324;
      end
    end else begin
      plru2_44 <= _GEN_876;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_45 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_45 <= _GEN_877;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_45 <= _GEN_877;
      end else begin
        plru2_45 <= _GEN_1325;
      end
    end else begin
      plru2_45 <= _GEN_877;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_46 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_46 <= _GEN_878;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_46 <= _GEN_878;
      end else begin
        plru2_46 <= _GEN_1326;
      end
    end else begin
      plru2_46 <= _GEN_878;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_47 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_47 <= _GEN_879;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_47 <= _GEN_879;
      end else begin
        plru2_47 <= _GEN_1327;
      end
    end else begin
      plru2_47 <= _GEN_879;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_48 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_48 <= _GEN_880;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_48 <= _GEN_880;
      end else begin
        plru2_48 <= _GEN_1328;
      end
    end else begin
      plru2_48 <= _GEN_880;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_49 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_49 <= _GEN_881;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_49 <= _GEN_881;
      end else begin
        plru2_49 <= _GEN_1329;
      end
    end else begin
      plru2_49 <= _GEN_881;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_50 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_50 <= _GEN_882;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_50 <= _GEN_882;
      end else begin
        plru2_50 <= _GEN_1330;
      end
    end else begin
      plru2_50 <= _GEN_882;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_51 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_51 <= _GEN_883;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_51 <= _GEN_883;
      end else begin
        plru2_51 <= _GEN_1331;
      end
    end else begin
      plru2_51 <= _GEN_883;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_52 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_52 <= _GEN_884;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_52 <= _GEN_884;
      end else begin
        plru2_52 <= _GEN_1332;
      end
    end else begin
      plru2_52 <= _GEN_884;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_53 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_53 <= _GEN_885;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_53 <= _GEN_885;
      end else begin
        plru2_53 <= _GEN_1333;
      end
    end else begin
      plru2_53 <= _GEN_885;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_54 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_54 <= _GEN_886;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_54 <= _GEN_886;
      end else begin
        plru2_54 <= _GEN_1334;
      end
    end else begin
      plru2_54 <= _GEN_886;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_55 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_55 <= _GEN_887;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_55 <= _GEN_887;
      end else begin
        plru2_55 <= _GEN_1335;
      end
    end else begin
      plru2_55 <= _GEN_887;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_56 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_56 <= _GEN_888;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_56 <= _GEN_888;
      end else begin
        plru2_56 <= _GEN_1336;
      end
    end else begin
      plru2_56 <= _GEN_888;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_57 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_57 <= _GEN_889;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_57 <= _GEN_889;
      end else begin
        plru2_57 <= _GEN_1337;
      end
    end else begin
      plru2_57 <= _GEN_889;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_58 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_58 <= _GEN_890;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_58 <= _GEN_890;
      end else begin
        plru2_58 <= _GEN_1338;
      end
    end else begin
      plru2_58 <= _GEN_890;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_59 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_59 <= _GEN_891;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_59 <= _GEN_891;
      end else begin
        plru2_59 <= _GEN_1339;
      end
    end else begin
      plru2_59 <= _GEN_891;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_60 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_60 <= _GEN_892;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_60 <= _GEN_892;
      end else begin
        plru2_60 <= _GEN_1340;
      end
    end else begin
      plru2_60 <= _GEN_892;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_61 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_61 <= _GEN_893;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_61 <= _GEN_893;
      end else begin
        plru2_61 <= _GEN_1341;
      end
    end else begin
      plru2_61 <= _GEN_893;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_62 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_62 <= _GEN_894;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_62 <= _GEN_894;
      end else begin
        plru2_62 <= _GEN_1342;
      end
    end else begin
      plru2_62 <= _GEN_894;
    end
    if (reset) begin // @[Cache_Soc.scala 91:22]
      plru2_63 <= 1'h0; // @[Cache_Soc.scala 91:22]
    end else if (state == 3'h4 & io_out_ret_valid & _cache_hit_T_2) begin // @[Cache_Soc.scala 106:61]
      if (_plru0_T_1) begin // @[Cache_Soc.scala 108:32]
        plru2_63 <= _GEN_895;
      end else if (_plru0_T_2) begin // @[Cache_Soc.scala 110:39]
        plru2_63 <= _GEN_895;
      end else begin
        plru2_63 <= _GEN_1343;
      end
    end else begin
      plru2_63 <= _GEN_895;
    end
    if (reset) begin // @[Cache_Soc.scala 296:24]
      counter <= 8'h0; // @[Cache_Soc.scala 296:24]
    end else if (!(_T_73)) begin // @[Conditional.scala 40:58]
      if (!(_T_74)) begin // @[Conditional.scala 39:67]
        if (_T_78) begin // @[Conditional.scala 39:67]
          counter <= _GEN_2351;
        end else begin
          counter <= _GEN_2374;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  wb_state = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  fence_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  rb_op = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  rb_uncache = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  rb_index = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  rb_tag = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  rb_offset = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  rb_wstrb = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  rb_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  wb_hitway = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  wb_index = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  wb_offset = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  wb_wstrb = _RAND_13[7:0];
  _RAND_14 = {2{`RANDOM}};
  wb_wdata = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  replace_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  replace_dirty = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  replace_tag = _RAND_17[21:0];
  _RAND_18 = {4{`RANDOM}};
  replace_data = _RAND_18[127:0];
  _RAND_19 = {1{`RANDOM}};
  plru0_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  plru0_1 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  plru0_2 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  plru0_3 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  plru0_4 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  plru0_5 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  plru0_6 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  plru0_7 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  plru0_8 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  plru0_9 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  plru0_10 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  plru0_11 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  plru0_12 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  plru0_13 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  plru0_14 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  plru0_15 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  plru0_16 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  plru0_17 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  plru0_18 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  plru0_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  plru0_20 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  plru0_21 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  plru0_22 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  plru0_23 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  plru0_24 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  plru0_25 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  plru0_26 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  plru0_27 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  plru0_28 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  plru0_29 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  plru0_30 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  plru0_31 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  plru0_32 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  plru0_33 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  plru0_34 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  plru0_35 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  plru0_36 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  plru0_37 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  plru0_38 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  plru0_39 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  plru0_40 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  plru0_41 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  plru0_42 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  plru0_43 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  plru0_44 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  plru0_45 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  plru0_46 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  plru0_47 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  plru0_48 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  plru0_49 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  plru0_50 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  plru0_51 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  plru0_52 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  plru0_53 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  plru0_54 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  plru0_55 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  plru0_56 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  plru0_57 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  plru0_58 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  plru0_59 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  plru0_60 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  plru0_61 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  plru0_62 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  plru0_63 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  plru1_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  plru1_1 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  plru1_2 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  plru1_3 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  plru1_4 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  plru1_5 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  plru1_6 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  plru1_7 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  plru1_8 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  plru1_9 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  plru1_10 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  plru1_11 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  plru1_12 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  plru1_13 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  plru1_14 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  plru1_15 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  plru1_16 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  plru1_17 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  plru1_18 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  plru1_19 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  plru1_20 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  plru1_21 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  plru1_22 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  plru1_23 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  plru1_24 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  plru1_25 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  plru1_26 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  plru1_27 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  plru1_28 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  plru1_29 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  plru1_30 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  plru1_31 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  plru1_32 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  plru1_33 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  plru1_34 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  plru1_35 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  plru1_36 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  plru1_37 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  plru1_38 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  plru1_39 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  plru1_40 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  plru1_41 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  plru1_42 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  plru1_43 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  plru1_44 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  plru1_45 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  plru1_46 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  plru1_47 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  plru1_48 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  plru1_49 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  plru1_50 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  plru1_51 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  plru1_52 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  plru1_53 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  plru1_54 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  plru1_55 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  plru1_56 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  plru1_57 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  plru1_58 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  plru1_59 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  plru1_60 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  plru1_61 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  plru1_62 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  plru1_63 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  plru2_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  plru2_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  plru2_2 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  plru2_3 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  plru2_4 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  plru2_5 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  plru2_6 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  plru2_7 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  plru2_8 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  plru2_9 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  plru2_10 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  plru2_11 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  plru2_12 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  plru2_13 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  plru2_14 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  plru2_15 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  plru2_16 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  plru2_17 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  plru2_18 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  plru2_19 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  plru2_20 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  plru2_21 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  plru2_22 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  plru2_23 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  plru2_24 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  plru2_25 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  plru2_26 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  plru2_27 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  plru2_28 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  plru2_29 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  plru2_30 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  plru2_31 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  plru2_32 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  plru2_33 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  plru2_34 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  plru2_35 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  plru2_36 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  plru2_37 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  plru2_38 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  plru2_39 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  plru2_40 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  plru2_41 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  plru2_42 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  plru2_43 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  plru2_44 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  plru2_45 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  plru2_46 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  plru2_47 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  plru2_48 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  plru2_49 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  plru2_50 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  plru2_51 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  plru2_52 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  plru2_53 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  plru2_54 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  plru2_55 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  plru2_56 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  plru2_57 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  plru2_58 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  plru2_59 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  plru2_60 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  plru2_61 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  plru2_62 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  plru2_63 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  counter = _RAND_211[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core_Soc(
  input          clock,
  input          reset,
  output         io_icache_bridge_rd_req,
  output [2:0]   io_icache_bridge_rd_size,
  output [31:0]  io_icache_bridge_rd_addr,
  input          io_icache_bridge_rd_rdy,
  input          io_icache_bridge_ret_valid,
  input  [127:0] io_icache_bridge_ret_data,
  output         io_dcache_bridge_rd_req,
  output [2:0]   io_dcache_bridge_rd_size,
  output [31:0]  io_dcache_bridge_rd_addr,
  input          io_dcache_bridge_rd_rdy,
  input          io_dcache_bridge_ret_valid,
  input  [127:0] io_dcache_bridge_ret_data,
  output         io_dcache_bridge_wr_req,
  output [2:0]   io_dcache_bridge_wr_size,
  output [31:0]  io_dcache_bridge_wr_addr,
  output [7:0]   io_dcache_bridge_wr_wstrb,
  output [127:0] io_dcache_bridge_wr_data,
  input          io_dcache_bridge_wr_rdy,
  input          io_dcache_bridge_wr_ok,
  output         io_sram_0_en,
  output         io_sram_0_wen,
  output [5:0]   io_sram_0_addr,
  output [127:0] io_sram_0_wdata,
  input  [127:0] io_sram_0_rdata,
  output         io_sram_1_en,
  output         io_sram_1_wen,
  output [5:0]   io_sram_1_addr,
  output [127:0] io_sram_1_wdata,
  input  [127:0] io_sram_1_rdata,
  output         io_sram_2_en,
  output         io_sram_2_wen,
  output [5:0]   io_sram_2_addr,
  output [127:0] io_sram_2_wdata,
  input  [127:0] io_sram_2_rdata,
  output         io_sram_3_en,
  output         io_sram_3_wen,
  output [5:0]   io_sram_3_addr,
  output [127:0] io_sram_3_wdata,
  input  [127:0] io_sram_3_rdata,
  output         io_sram_4_en,
  output         io_sram_4_wen,
  output [5:0]   io_sram_4_addr,
  output [127:0] io_sram_4_wdata,
  input  [127:0] io_sram_4_rdata,
  output         io_sram_5_en,
  output         io_sram_5_wen,
  output [5:0]   io_sram_5_addr,
  output [127:0] io_sram_5_wdata,
  input  [127:0] io_sram_5_rdata,
  output         io_sram_6_en,
  output         io_sram_6_wen,
  output [5:0]   io_sram_6_addr,
  output [127:0] io_sram_6_wdata,
  input  [127:0] io_sram_6_rdata,
  output         io_sram_7_en,
  output         io_sram_7_wen,
  output [5:0]   io_sram_7_addr,
  output [127:0] io_sram_7_wdata,
  input  [127:0] io_sram_7_rdata,
  output [31:0]  io_commit_0_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[Core.scala 12:19]
  wire  ifu_reset; // @[Core.scala 12:19]
  wire  ifu_io_imem_valid; // @[Core.scala 12:19]
  wire [31:0] ifu_io_imem_addr; // @[Core.scala 12:19]
  wire  ifu_io_imem_fence; // @[Core.scala 12:19]
  wire  ifu_io_imem_fence_finish; // @[Core.scala 12:19]
  wire  ifu_io_imem_data_ok; // @[Core.scala 12:19]
  wire [127:0] ifu_io_imem_inst; // @[Core.scala 12:19]
  wire  ifu_io_out_ready; // @[Core.scala 12:19]
  wire  ifu_io_out_valid; // @[Core.scala 12:19]
  wire [31:0] ifu_io_out_bits_pc; // @[Core.scala 12:19]
  wire [127:0] ifu_io_out_bits_inst; // @[Core.scala 12:19]
  wire  ifu_io_out_bits_uncache; // @[Core.scala 12:19]
  wire [1:0] ifu_io_out_bits_offset; // @[Core.scala 12:19]
  wire [1:0] ifu_io_out_bits_bp_br_offset; // @[Core.scala 12:19]
  wire  ifu_io_out_bits_bp_br_taken; // @[Core.scala 12:19]
  wire [31:0] ifu_io_out_bits_bp_br_target; // @[Core.scala 12:19]
  wire [1:0] ifu_io_out_bits_bp_br_type; // @[Core.scala 12:19]
  wire  ifu_io_reflush_bus_is_reflush; // @[Core.scala 12:19]
  wire [31:0] ifu_io_reflush_bus_br_target; // @[Core.scala 12:19]
  wire  ifu_io_bpu_valid; // @[Core.scala 12:19]
  wire [31:0] ifu_io_bpu_pc; // @[Core.scala 12:19]
  wire  ifu_io_bpu_bp_ok; // @[Core.scala 12:19]
  wire  ifu_io_bpu_bp_taken; // @[Core.scala 12:19]
  wire [31:0] ifu_io_bpu_bp_target; // @[Core.scala 12:19]
  wire [1:0] ifu_io_bpu_bp_offset; // @[Core.scala 12:19]
  wire  ifu_io_bpu_is_reflush; // @[Core.scala 12:19]
  wire [1:0] ifu_io_bpu_bp_type; // @[Core.scala 12:19]
  wire [2:0] ifu_io_bpu_call_count; // @[Core.scala 12:19]
  wire [2:0] ifu_io_bpu_ret_count; // @[Core.scala 12:19]
  wire  ifu_dcache_fence_finish_0; // @[Core.scala 12:19]
  wire  ifu_fence_i; // @[Core.scala 12:19]
  wire  ifu_icache_fence_finish_0; // @[Core.scala 12:19]
  wire  iqueue_clock; // @[Core.scala 13:22]
  wire  iqueue_reset; // @[Core.scala 13:22]
  wire  iqueue_io_in_ready; // @[Core.scala 13:22]
  wire  iqueue_io_in_valid; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_in_bits_pc; // @[Core.scala 13:22]
  wire [127:0] iqueue_io_in_bits_inst; // @[Core.scala 13:22]
  wire  iqueue_io_in_bits_uncache; // @[Core.scala 13:22]
  wire [1:0] iqueue_io_in_bits_offset; // @[Core.scala 13:22]
  wire [1:0] iqueue_io_in_bits_bp_br_offset; // @[Core.scala 13:22]
  wire  iqueue_io_in_bits_bp_br_taken; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_in_bits_bp_br_target; // @[Core.scala 13:22]
  wire [1:0] iqueue_io_in_bits_bp_br_type; // @[Core.scala 13:22]
  wire  iqueue_io_out_ready; // @[Core.scala 13:22]
  wire  iqueue_io_out_valid; // @[Core.scala 13:22]
  wire  iqueue_io_out_bits_0_valid; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_out_bits_0_pc; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_out_bits_0_inst; // @[Core.scala 13:22]
  wire  iqueue_io_out_bits_0_bp_br_taken; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_out_bits_0_bp_br_target; // @[Core.scala 13:22]
  wire [1:0] iqueue_io_out_bits_0_bp_br_type; // @[Core.scala 13:22]
  wire  iqueue_io_out_bits_1_valid; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_out_bits_1_pc; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_out_bits_1_inst; // @[Core.scala 13:22]
  wire  iqueue_io_out_bits_1_bp_br_taken; // @[Core.scala 13:22]
  wire [31:0] iqueue_io_out_bits_1_bp_br_target; // @[Core.scala 13:22]
  wire [1:0] iqueue_io_out_bits_1_bp_br_type; // @[Core.scala 13:22]
  wire  iqueue_frontend_reflush; // @[Core.scala 13:22]
  wire  idu_clock; // @[Core.scala 14:19]
  wire  idu_reset; // @[Core.scala 14:19]
  wire  idu_io_in_ready; // @[Core.scala 14:19]
  wire  idu_io_in_valid; // @[Core.scala 14:19]
  wire  idu_io_in_bits_0_valid; // @[Core.scala 14:19]
  wire [31:0] idu_io_in_bits_0_pc; // @[Core.scala 14:19]
  wire [31:0] idu_io_in_bits_0_inst; // @[Core.scala 14:19]
  wire  idu_io_in_bits_0_bp_br_taken; // @[Core.scala 14:19]
  wire [31:0] idu_io_in_bits_0_bp_br_target; // @[Core.scala 14:19]
  wire [1:0] idu_io_in_bits_0_bp_br_type; // @[Core.scala 14:19]
  wire  idu_io_in_bits_1_valid; // @[Core.scala 14:19]
  wire [31:0] idu_io_in_bits_1_pc; // @[Core.scala 14:19]
  wire [31:0] idu_io_in_bits_1_inst; // @[Core.scala 14:19]
  wire  idu_io_in_bits_1_bp_br_taken; // @[Core.scala 14:19]
  wire [31:0] idu_io_in_bits_1_bp_br_target; // @[Core.scala 14:19]
  wire [1:0] idu_io_in_bits_1_bp_br_type; // @[Core.scala 14:19]
  wire  idu_io_out_ready; // @[Core.scala 14:19]
  wire  idu_io_out_valid; // @[Core.scala 14:19]
  wire  idu_io_out_bits_0_valid; // @[Core.scala 14:19]
  wire [31:0] idu_io_out_bits_0_pc; // @[Core.scala 14:19]
  wire [31:0] idu_io_out_bits_0_inst; // @[Core.scala 14:19]
  wire [1:0] idu_io_out_bits_0_src1; // @[Core.scala 14:19]
  wire [1:0] idu_io_out_bits_0_src2; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_0_rs1; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_0_rs2; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_0_dest; // @[Core.scala 14:19]
  wire [63:0] idu_io_out_bits_0_imm; // @[Core.scala 14:19]
  wire [2:0] idu_io_out_bits_0_fu_type; // @[Core.scala 14:19]
  wire [3:0] idu_io_out_bits_0_bru_op; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_0_alu_op; // @[Core.scala 14:19]
  wire [3:0] idu_io_out_bits_0_lsu_op; // @[Core.scala 14:19]
  wire [2:0] idu_io_out_bits_0_csr_op; // @[Core.scala 14:19]
  wire [3:0] idu_io_out_bits_0_mdu_op; // @[Core.scala 14:19]
  wire  idu_io_out_bits_0_wen; // @[Core.scala 14:19]
  wire  idu_io_out_bits_0_rv64; // @[Core.scala 14:19]
  wire  idu_io_out_bits_0_bp_br_taken; // @[Core.scala 14:19]
  wire [31:0] idu_io_out_bits_0_bp_br_target; // @[Core.scala 14:19]
  wire [1:0] idu_io_out_bits_0_bp_br_type; // @[Core.scala 14:19]
  wire  idu_io_out_bits_1_valid; // @[Core.scala 14:19]
  wire [31:0] idu_io_out_bits_1_pc; // @[Core.scala 14:19]
  wire [31:0] idu_io_out_bits_1_inst; // @[Core.scala 14:19]
  wire [1:0] idu_io_out_bits_1_src1; // @[Core.scala 14:19]
  wire [1:0] idu_io_out_bits_1_src2; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_1_rs1; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_1_rs2; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_1_dest; // @[Core.scala 14:19]
  wire [63:0] idu_io_out_bits_1_imm; // @[Core.scala 14:19]
  wire [2:0] idu_io_out_bits_1_fu_type; // @[Core.scala 14:19]
  wire [3:0] idu_io_out_bits_1_bru_op; // @[Core.scala 14:19]
  wire [4:0] idu_io_out_bits_1_alu_op; // @[Core.scala 14:19]
  wire [3:0] idu_io_out_bits_1_lsu_op; // @[Core.scala 14:19]
  wire [2:0] idu_io_out_bits_1_csr_op; // @[Core.scala 14:19]
  wire [3:0] idu_io_out_bits_1_mdu_op; // @[Core.scala 14:19]
  wire  idu_io_out_bits_1_wen; // @[Core.scala 14:19]
  wire  idu_io_out_bits_1_rv64; // @[Core.scala 14:19]
  wire  idu_io_out_bits_1_bp_br_taken; // @[Core.scala 14:19]
  wire [31:0] idu_io_out_bits_1_bp_br_target; // @[Core.scala 14:19]
  wire [1:0] idu_io_out_bits_1_bp_br_type; // @[Core.scala 14:19]
  wire  idu_frontend_reflush; // @[Core.scala 14:19]
  wire  issue_clock; // @[Core.scala 15:21]
  wire  issue_reset; // @[Core.scala 15:21]
  wire  issue_io_in_ready; // @[Core.scala 15:21]
  wire  issue_io_in_valid; // @[Core.scala 15:21]
  wire  issue_io_in_bits_0_valid; // @[Core.scala 15:21]
  wire [31:0] issue_io_in_bits_0_pc; // @[Core.scala 15:21]
  wire [31:0] issue_io_in_bits_0_inst; // @[Core.scala 15:21]
  wire [1:0] issue_io_in_bits_0_src1; // @[Core.scala 15:21]
  wire [1:0] issue_io_in_bits_0_src2; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_0_rs1; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_0_rs2; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_0_dest; // @[Core.scala 15:21]
  wire [63:0] issue_io_in_bits_0_imm; // @[Core.scala 15:21]
  wire [2:0] issue_io_in_bits_0_fu_type; // @[Core.scala 15:21]
  wire [3:0] issue_io_in_bits_0_bru_op; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_0_alu_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_in_bits_0_lsu_op; // @[Core.scala 15:21]
  wire [2:0] issue_io_in_bits_0_csr_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_in_bits_0_mdu_op; // @[Core.scala 15:21]
  wire  issue_io_in_bits_0_wen; // @[Core.scala 15:21]
  wire  issue_io_in_bits_0_rv64; // @[Core.scala 15:21]
  wire  issue_io_in_bits_0_bp_br_taken; // @[Core.scala 15:21]
  wire [31:0] issue_io_in_bits_0_bp_br_target; // @[Core.scala 15:21]
  wire [1:0] issue_io_in_bits_0_bp_br_type; // @[Core.scala 15:21]
  wire  issue_io_in_bits_1_valid; // @[Core.scala 15:21]
  wire [31:0] issue_io_in_bits_1_pc; // @[Core.scala 15:21]
  wire [31:0] issue_io_in_bits_1_inst; // @[Core.scala 15:21]
  wire [1:0] issue_io_in_bits_1_src1; // @[Core.scala 15:21]
  wire [1:0] issue_io_in_bits_1_src2; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_1_rs1; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_1_rs2; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_1_dest; // @[Core.scala 15:21]
  wire [63:0] issue_io_in_bits_1_imm; // @[Core.scala 15:21]
  wire [2:0] issue_io_in_bits_1_fu_type; // @[Core.scala 15:21]
  wire [3:0] issue_io_in_bits_1_bru_op; // @[Core.scala 15:21]
  wire [4:0] issue_io_in_bits_1_alu_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_in_bits_1_lsu_op; // @[Core.scala 15:21]
  wire [2:0] issue_io_in_bits_1_csr_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_in_bits_1_mdu_op; // @[Core.scala 15:21]
  wire  issue_io_in_bits_1_wen; // @[Core.scala 15:21]
  wire  issue_io_in_bits_1_rv64; // @[Core.scala 15:21]
  wire  issue_io_in_bits_1_bp_br_taken; // @[Core.scala 15:21]
  wire [31:0] issue_io_in_bits_1_bp_br_target; // @[Core.scala 15:21]
  wire [1:0] issue_io_in_bits_1_bp_br_type; // @[Core.scala 15:21]
  wire  issue_io_out_ready; // @[Core.scala 15:21]
  wire  issue_io_out_valid; // @[Core.scala 15:21]
  wire  issue_io_out_bits_0_valid; // @[Core.scala 15:21]
  wire [31:0] issue_io_out_bits_0_pc; // @[Core.scala 15:21]
  wire [31:0] issue_io_out_bits_0_inst; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_0_src1_value; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_0_src2_value; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_0_rs2_value; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_0_imm; // @[Core.scala 15:21]
  wire [4:0] issue_io_out_bits_0_rs1; // @[Core.scala 15:21]
  wire [4:0] issue_io_out_bits_0_dest; // @[Core.scala 15:21]
  wire [2:0] issue_io_out_bits_0_fu_type; // @[Core.scala 15:21]
  wire [3:0] issue_io_out_bits_0_bru_op; // @[Core.scala 15:21]
  wire [4:0] issue_io_out_bits_0_alu_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_out_bits_0_lsu_op; // @[Core.scala 15:21]
  wire [2:0] issue_io_out_bits_0_csr_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_out_bits_0_mdu_op; // @[Core.scala 15:21]
  wire  issue_io_out_bits_0_wen; // @[Core.scala 15:21]
  wire  issue_io_out_bits_0_rv64; // @[Core.scala 15:21]
  wire  issue_io_out_bits_0_bp_br_taken; // @[Core.scala 15:21]
  wire [31:0] issue_io_out_bits_0_bp_br_target; // @[Core.scala 15:21]
  wire [1:0] issue_io_out_bits_0_bp_br_type; // @[Core.scala 15:21]
  wire  issue_io_out_bits_1_valid; // @[Core.scala 15:21]
  wire [31:0] issue_io_out_bits_1_pc; // @[Core.scala 15:21]
  wire [31:0] issue_io_out_bits_1_inst; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_1_src1_value; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_1_src2_value; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_1_rs2_value; // @[Core.scala 15:21]
  wire [63:0] issue_io_out_bits_1_imm; // @[Core.scala 15:21]
  wire [4:0] issue_io_out_bits_1_rs1; // @[Core.scala 15:21]
  wire [4:0] issue_io_out_bits_1_dest; // @[Core.scala 15:21]
  wire [2:0] issue_io_out_bits_1_fu_type; // @[Core.scala 15:21]
  wire [3:0] issue_io_out_bits_1_bru_op; // @[Core.scala 15:21]
  wire [4:0] issue_io_out_bits_1_alu_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_out_bits_1_lsu_op; // @[Core.scala 15:21]
  wire [2:0] issue_io_out_bits_1_csr_op; // @[Core.scala 15:21]
  wire [3:0] issue_io_out_bits_1_mdu_op; // @[Core.scala 15:21]
  wire  issue_io_out_bits_1_wen; // @[Core.scala 15:21]
  wire  issue_io_out_bits_1_rv64; // @[Core.scala 15:21]
  wire  issue_io_out_bits_1_bp_br_taken; // @[Core.scala 15:21]
  wire [31:0] issue_io_out_bits_1_bp_br_target; // @[Core.scala 15:21]
  wire [1:0] issue_io_out_bits_1_bp_br_type; // @[Core.scala 15:21]
  wire  issue_io_wb_bus_0_rf_wen; // @[Core.scala 15:21]
  wire [4:0] issue_io_wb_bus_0_rf_waddr; // @[Core.scala 15:21]
  wire [63:0] issue_io_wb_bus_0_rf_wdata; // @[Core.scala 15:21]
  wire  issue_io_wb_bus_1_rf_wen; // @[Core.scala 15:21]
  wire [4:0] issue_io_wb_bus_1_rf_waddr; // @[Core.scala 15:21]
  wire [63:0] issue_io_wb_bus_1_rf_wdata; // @[Core.scala 15:21]
  wire  issue_io_ex_fwd_0_blk_valid; // @[Core.scala 15:21]
  wire  issue_io_ex_fwd_0_fwd_valid; // @[Core.scala 15:21]
  wire [4:0] issue_io_ex_fwd_0_rf_waddr; // @[Core.scala 15:21]
  wire [63:0] issue_io_ex_fwd_0_rf_wdata; // @[Core.scala 15:21]
  wire  issue_io_ex_fwd_1_blk_valid; // @[Core.scala 15:21]
  wire  issue_io_ex_fwd_1_fwd_valid; // @[Core.scala 15:21]
  wire [4:0] issue_io_ex_fwd_1_rf_waddr; // @[Core.scala 15:21]
  wire [63:0] issue_io_ex_fwd_1_rf_wdata; // @[Core.scala 15:21]
  wire  issue_frontend_reflush; // @[Core.scala 15:21]
  wire  exu_clock; // @[Core.scala 16:19]
  wire  exu_reset; // @[Core.scala 16:19]
  wire  exu_io_dmem_valid; // @[Core.scala 16:19]
  wire  exu_io_dmem_op; // @[Core.scala 16:19]
  wire [31:0] exu_io_dmem_addr; // @[Core.scala 16:19]
  wire [7:0] exu_io_dmem_wstrb; // @[Core.scala 16:19]
  wire [63:0] exu_io_dmem_wdata; // @[Core.scala 16:19]
  wire  exu_io_dmem_fence; // @[Core.scala 16:19]
  wire  exu_io_dmem_fence_finish; // @[Core.scala 16:19]
  wire  exu_io_dmem_data_ok; // @[Core.scala 16:19]
  wire [63:0] exu_io_dmem_rdata; // @[Core.scala 16:19]
  wire  exu_io_in_ready; // @[Core.scala 16:19]
  wire  exu_io_in_valid; // @[Core.scala 16:19]
  wire  exu_io_in_bits_0_valid; // @[Core.scala 16:19]
  wire [31:0] exu_io_in_bits_0_pc; // @[Core.scala 16:19]
  wire [31:0] exu_io_in_bits_0_inst; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_0_src1_value; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_0_src2_value; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_0_rs2_value; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_0_imm; // @[Core.scala 16:19]
  wire [4:0] exu_io_in_bits_0_rs1; // @[Core.scala 16:19]
  wire [4:0] exu_io_in_bits_0_dest; // @[Core.scala 16:19]
  wire [2:0] exu_io_in_bits_0_fu_type; // @[Core.scala 16:19]
  wire [3:0] exu_io_in_bits_0_bru_op; // @[Core.scala 16:19]
  wire [4:0] exu_io_in_bits_0_alu_op; // @[Core.scala 16:19]
  wire [3:0] exu_io_in_bits_0_lsu_op; // @[Core.scala 16:19]
  wire [2:0] exu_io_in_bits_0_csr_op; // @[Core.scala 16:19]
  wire [3:0] exu_io_in_bits_0_mdu_op; // @[Core.scala 16:19]
  wire  exu_io_in_bits_0_wen; // @[Core.scala 16:19]
  wire  exu_io_in_bits_0_rv64; // @[Core.scala 16:19]
  wire  exu_io_in_bits_0_bp_br_taken; // @[Core.scala 16:19]
  wire [31:0] exu_io_in_bits_0_bp_br_target; // @[Core.scala 16:19]
  wire [1:0] exu_io_in_bits_0_bp_br_type; // @[Core.scala 16:19]
  wire  exu_io_in_bits_1_valid; // @[Core.scala 16:19]
  wire [31:0] exu_io_in_bits_1_pc; // @[Core.scala 16:19]
  wire [31:0] exu_io_in_bits_1_inst; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_1_src1_value; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_1_src2_value; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_1_rs2_value; // @[Core.scala 16:19]
  wire [63:0] exu_io_in_bits_1_imm; // @[Core.scala 16:19]
  wire [4:0] exu_io_in_bits_1_rs1; // @[Core.scala 16:19]
  wire [4:0] exu_io_in_bits_1_dest; // @[Core.scala 16:19]
  wire [2:0] exu_io_in_bits_1_fu_type; // @[Core.scala 16:19]
  wire [3:0] exu_io_in_bits_1_bru_op; // @[Core.scala 16:19]
  wire [4:0] exu_io_in_bits_1_alu_op; // @[Core.scala 16:19]
  wire [3:0] exu_io_in_bits_1_lsu_op; // @[Core.scala 16:19]
  wire [2:0] exu_io_in_bits_1_csr_op; // @[Core.scala 16:19]
  wire [3:0] exu_io_in_bits_1_mdu_op; // @[Core.scala 16:19]
  wire  exu_io_in_bits_1_wen; // @[Core.scala 16:19]
  wire  exu_io_in_bits_1_rv64; // @[Core.scala 16:19]
  wire  exu_io_in_bits_1_bp_br_taken; // @[Core.scala 16:19]
  wire [31:0] exu_io_in_bits_1_bp_br_target; // @[Core.scala 16:19]
  wire [1:0] exu_io_in_bits_1_bp_br_type; // @[Core.scala 16:19]
  wire  exu_io_out_valid; // @[Core.scala 16:19]
  wire  exu_io_out_bits_0_valid; // @[Core.scala 16:19]
  wire [31:0] exu_io_out_bits_0_pc; // @[Core.scala 16:19]
  wire [63:0] exu_io_out_bits_0_final_result; // @[Core.scala 16:19]
  wire [4:0] exu_io_out_bits_0_dest; // @[Core.scala 16:19]
  wire  exu_io_out_bits_0_wen; // @[Core.scala 16:19]
  wire  exu_io_out_bits_1_valid; // @[Core.scala 16:19]
  wire [63:0] exu_io_out_bits_1_final_result; // @[Core.scala 16:19]
  wire [4:0] exu_io_out_bits_1_dest; // @[Core.scala 16:19]
  wire  exu_io_out_bits_1_wen; // @[Core.scala 16:19]
  wire  exu_io_forward_0_blk_valid; // @[Core.scala 16:19]
  wire  exu_io_forward_0_fwd_valid; // @[Core.scala 16:19]
  wire [4:0] exu_io_forward_0_rf_waddr; // @[Core.scala 16:19]
  wire [63:0] exu_io_forward_0_rf_wdata; // @[Core.scala 16:19]
  wire  exu_io_forward_1_blk_valid; // @[Core.scala 16:19]
  wire  exu_io_forward_1_fwd_valid; // @[Core.scala 16:19]
  wire [4:0] exu_io_forward_1_rf_waddr; // @[Core.scala 16:19]
  wire [63:0] exu_io_forward_1_rf_wdata; // @[Core.scala 16:19]
  wire  exu_io_reflush_bus_is_reflush; // @[Core.scala 16:19]
  wire [31:0] exu_io_reflush_bus_br_target; // @[Core.scala 16:19]
  wire  exu_io_bpu_valid; // @[Core.scala 16:19]
  wire [31:0] exu_io_bpu_pc; // @[Core.scala 16:19]
  wire  exu_io_bpu_bp_taken; // @[Core.scala 16:19]
  wire [31:0] exu_io_bpu_bp_target; // @[Core.scala 16:19]
  wire [1:0] exu_io_bpu_bp_type; // @[Core.scala 16:19]
  wire  exu_io_bpu_bp_wrong; // @[Core.scala 16:19]
  wire  exu_io_bpu_fence; // @[Core.scala 16:19]
  wire [2:0] exu_io_bpu_call_count; // @[Core.scala 16:19]
  wire [2:0] exu_io_bpu_ret_count; // @[Core.scala 16:19]
  wire  exu_frontend_reflush_0; // @[Core.scala 16:19]
  wire  exu_dcache_fence_finish; // @[Core.scala 16:19]
  wire  exu_fence_0; // @[Core.scala 16:19]
  wire  exu_icache_fence_finish; // @[Core.scala 16:19]
  wire  wbu_io__in_valid; // @[Core.scala 17:19]
  wire  wbu_io__in_bits_0_valid; // @[Core.scala 17:19]
  wire [31:0] wbu_io__in_bits_0_pc; // @[Core.scala 17:19]
  wire [63:0] wbu_io__in_bits_0_final_result; // @[Core.scala 17:19]
  wire [4:0] wbu_io__in_bits_0_dest; // @[Core.scala 17:19]
  wire  wbu_io__in_bits_0_wen; // @[Core.scala 17:19]
  wire  wbu_io__in_bits_1_valid; // @[Core.scala 17:19]
  wire [63:0] wbu_io__in_bits_1_final_result; // @[Core.scala 17:19]
  wire [4:0] wbu_io__in_bits_1_dest; // @[Core.scala 17:19]
  wire  wbu_io__in_bits_1_wen; // @[Core.scala 17:19]
  wire  wbu_io__wb_bus_0_rf_wen; // @[Core.scala 17:19]
  wire [4:0] wbu_io__wb_bus_0_rf_waddr; // @[Core.scala 17:19]
  wire [63:0] wbu_io__wb_bus_0_rf_wdata; // @[Core.scala 17:19]
  wire  wbu_io__wb_bus_1_rf_wen; // @[Core.scala 17:19]
  wire [4:0] wbu_io__wb_bus_1_rf_waddr; // @[Core.scala 17:19]
  wire [63:0] wbu_io__wb_bus_1_rf_wdata; // @[Core.scala 17:19]
  wire [31:0] wbu_io__commit_0_pc; // @[Core.scala 17:19]
  wire [31:0] wbu_io_commit_0_pc; // @[Core.scala 17:19]
  wire  bpu_clock; // @[Core.scala 18:19]
  wire  bpu_reset; // @[Core.scala 18:19]
  wire  bpu_io_ifu_valid; // @[Core.scala 18:19]
  wire [31:0] bpu_io_ifu_pc; // @[Core.scala 18:19]
  wire  bpu_io_ifu_bp_ok; // @[Core.scala 18:19]
  wire  bpu_io_ifu_bp_taken; // @[Core.scala 18:19]
  wire [31:0] bpu_io_ifu_bp_target; // @[Core.scala 18:19]
  wire [1:0] bpu_io_ifu_bp_offset; // @[Core.scala 18:19]
  wire  bpu_io_ifu_is_reflush; // @[Core.scala 18:19]
  wire [1:0] bpu_io_ifu_bp_type; // @[Core.scala 18:19]
  wire [2:0] bpu_io_ifu_call_count; // @[Core.scala 18:19]
  wire [2:0] bpu_io_ifu_ret_count; // @[Core.scala 18:19]
  wire  bpu_io_exu_valid; // @[Core.scala 18:19]
  wire [31:0] bpu_io_exu_pc; // @[Core.scala 18:19]
  wire  bpu_io_exu_bp_taken; // @[Core.scala 18:19]
  wire [31:0] bpu_io_exu_bp_target; // @[Core.scala 18:19]
  wire [1:0] bpu_io_exu_bp_type; // @[Core.scala 18:19]
  wire  bpu_io_exu_bp_wrong; // @[Core.scala 18:19]
  wire  bpu_io_exu_fence; // @[Core.scala 18:19]
  wire [2:0] bpu_io_exu_call_count; // @[Core.scala 18:19]
  wire [2:0] bpu_io_exu_ret_count; // @[Core.scala 18:19]
  wire  icache_clock; // @[Core.scala 19:22]
  wire  icache_reset; // @[Core.scala 19:22]
  wire  icache_io_in_valid; // @[Core.scala 19:22]
  wire  icache_io_in_op; // @[Core.scala 19:22]
  wire [31:0] icache_io_in_addr; // @[Core.scala 19:22]
  wire [7:0] icache_io_in_wstrb; // @[Core.scala 19:22]
  wire [63:0] icache_io_in_wdata; // @[Core.scala 19:22]
  wire  icache_io_in_fence; // @[Core.scala 19:22]
  wire  icache_io_in_fence_finish; // @[Core.scala 19:22]
  wire  icache_io_in_data_ok; // @[Core.scala 19:22]
  wire [63:0] icache_io_in_rdata; // @[Core.scala 19:22]
  wire [127:0] icache_io_in_inst; // @[Core.scala 19:22]
  wire  icache_io_out_rd_req; // @[Core.scala 19:22]
  wire [2:0] icache_io_out_rd_size; // @[Core.scala 19:22]
  wire [31:0] icache_io_out_rd_addr; // @[Core.scala 19:22]
  wire  icache_io_out_rd_rdy; // @[Core.scala 19:22]
  wire  icache_io_out_ret_valid; // @[Core.scala 19:22]
  wire [127:0] icache_io_out_ret_data; // @[Core.scala 19:22]
  wire  icache_io_out_wr_req; // @[Core.scala 19:22]
  wire [2:0] icache_io_out_wr_size; // @[Core.scala 19:22]
  wire [31:0] icache_io_out_wr_addr; // @[Core.scala 19:22]
  wire [7:0] icache_io_out_wr_wstrb; // @[Core.scala 19:22]
  wire [127:0] icache_io_out_wr_data; // @[Core.scala 19:22]
  wire  icache_io_out_wr_rdy; // @[Core.scala 19:22]
  wire  icache_io_out_wr_ok; // @[Core.scala 19:22]
  wire  icache_io_sram_0_en; // @[Core.scala 19:22]
  wire  icache_io_sram_0_wen; // @[Core.scala 19:22]
  wire [5:0] icache_io_sram_0_addr; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_0_wdata; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_0_rdata; // @[Core.scala 19:22]
  wire  icache_io_sram_1_en; // @[Core.scala 19:22]
  wire  icache_io_sram_1_wen; // @[Core.scala 19:22]
  wire [5:0] icache_io_sram_1_addr; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_1_wdata; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_1_rdata; // @[Core.scala 19:22]
  wire  icache_io_sram_2_en; // @[Core.scala 19:22]
  wire  icache_io_sram_2_wen; // @[Core.scala 19:22]
  wire [5:0] icache_io_sram_2_addr; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_2_wdata; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_2_rdata; // @[Core.scala 19:22]
  wire  icache_io_sram_3_en; // @[Core.scala 19:22]
  wire  icache_io_sram_3_wen; // @[Core.scala 19:22]
  wire [5:0] icache_io_sram_3_addr; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_3_wdata; // @[Core.scala 19:22]
  wire [127:0] icache_io_sram_3_rdata; // @[Core.scala 19:22]
  wire  dcache_clock; // @[Core.scala 20:22]
  wire  dcache_reset; // @[Core.scala 20:22]
  wire  dcache_io_in_valid; // @[Core.scala 20:22]
  wire  dcache_io_in_op; // @[Core.scala 20:22]
  wire [31:0] dcache_io_in_addr; // @[Core.scala 20:22]
  wire [7:0] dcache_io_in_wstrb; // @[Core.scala 20:22]
  wire [63:0] dcache_io_in_wdata; // @[Core.scala 20:22]
  wire  dcache_io_in_fence; // @[Core.scala 20:22]
  wire  dcache_io_in_fence_finish; // @[Core.scala 20:22]
  wire  dcache_io_in_data_ok; // @[Core.scala 20:22]
  wire [63:0] dcache_io_in_rdata; // @[Core.scala 20:22]
  wire [127:0] dcache_io_in_inst; // @[Core.scala 20:22]
  wire  dcache_io_out_rd_req; // @[Core.scala 20:22]
  wire [2:0] dcache_io_out_rd_size; // @[Core.scala 20:22]
  wire [31:0] dcache_io_out_rd_addr; // @[Core.scala 20:22]
  wire  dcache_io_out_rd_rdy; // @[Core.scala 20:22]
  wire  dcache_io_out_ret_valid; // @[Core.scala 20:22]
  wire [127:0] dcache_io_out_ret_data; // @[Core.scala 20:22]
  wire  dcache_io_out_wr_req; // @[Core.scala 20:22]
  wire [2:0] dcache_io_out_wr_size; // @[Core.scala 20:22]
  wire [31:0] dcache_io_out_wr_addr; // @[Core.scala 20:22]
  wire [7:0] dcache_io_out_wr_wstrb; // @[Core.scala 20:22]
  wire [127:0] dcache_io_out_wr_data; // @[Core.scala 20:22]
  wire  dcache_io_out_wr_rdy; // @[Core.scala 20:22]
  wire  dcache_io_out_wr_ok; // @[Core.scala 20:22]
  wire  dcache_io_sram_0_en; // @[Core.scala 20:22]
  wire  dcache_io_sram_0_wen; // @[Core.scala 20:22]
  wire [5:0] dcache_io_sram_0_addr; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_0_wdata; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_0_rdata; // @[Core.scala 20:22]
  wire  dcache_io_sram_1_en; // @[Core.scala 20:22]
  wire  dcache_io_sram_1_wen; // @[Core.scala 20:22]
  wire [5:0] dcache_io_sram_1_addr; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_1_wdata; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_1_rdata; // @[Core.scala 20:22]
  wire  dcache_io_sram_2_en; // @[Core.scala 20:22]
  wire  dcache_io_sram_2_wen; // @[Core.scala 20:22]
  wire [5:0] dcache_io_sram_2_addr; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_2_wdata; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_2_rdata; // @[Core.scala 20:22]
  wire  dcache_io_sram_3_en; // @[Core.scala 20:22]
  wire  dcache_io_sram_3_wen; // @[Core.scala 20:22]
  wire [5:0] dcache_io_sram_3_addr; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_3_wdata; // @[Core.scala 20:22]
  wire [127:0] dcache_io_sram_3_rdata; // @[Core.scala 20:22]
  reg  valid; // @[Connect.scala 6:24]
  wire  fire = ifu_io_out_valid & iqueue_io_in_ready; // @[Connect.scala 7:27]
  wire  _T_1 = iqueue_io_in_ready & iqueue_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_0 = _T_1 ? 1'h0 : valid; // @[Connect.scala 8:23 Connect.scala 8:31 Connect.scala 6:24]
  wire  _GEN_1 = fire | _GEN_0; // @[Connect.scala 9:17 Connect.scala 9:25]
  wire  frontend_reflush_0 = exu_frontend_reflush_0;
  reg [31:0] iqueue_io_in_bits_r_pc; // @[Reg.scala 27:20]
  reg [127:0] iqueue_io_in_bits_r_inst; // @[Reg.scala 27:20]
  reg  iqueue_io_in_bits_r_uncache; // @[Reg.scala 27:20]
  reg [1:0] iqueue_io_in_bits_r_offset; // @[Reg.scala 27:20]
  reg [1:0] iqueue_io_in_bits_r_bp_br_offset; // @[Reg.scala 27:20]
  reg  iqueue_io_in_bits_r_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] iqueue_io_in_bits_r_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] iqueue_io_in_bits_r_bp_br_type; // @[Reg.scala 27:20]
  reg  valid_1; // @[Connect.scala 6:24]
  wire  fire_1 = iqueue_io_out_valid & idu_io_in_ready; // @[Connect.scala 7:27]
  wire  _T_3 = idu_io_in_ready & idu_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_11 = _T_3 ? 1'h0 : valid_1; // @[Connect.scala 8:23 Connect.scala 8:31 Connect.scala 6:24]
  wire  _GEN_12 = fire_1 | _GEN_11; // @[Connect.scala 9:17 Connect.scala 9:25]
  reg  idu_io_in_bits_r_0_valid; // @[Reg.scala 27:20]
  reg [31:0] idu_io_in_bits_r_0_pc; // @[Reg.scala 27:20]
  reg [31:0] idu_io_in_bits_r_0_inst; // @[Reg.scala 27:20]
  reg  idu_io_in_bits_r_0_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] idu_io_in_bits_r_0_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] idu_io_in_bits_r_0_bp_br_type; // @[Reg.scala 27:20]
  reg  idu_io_in_bits_r_1_valid; // @[Reg.scala 27:20]
  reg [31:0] idu_io_in_bits_r_1_pc; // @[Reg.scala 27:20]
  reg [31:0] idu_io_in_bits_r_1_inst; // @[Reg.scala 27:20]
  reg  idu_io_in_bits_r_1_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] idu_io_in_bits_r_1_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] idu_io_in_bits_r_1_bp_br_type; // @[Reg.scala 27:20]
  reg  valid_2; // @[Connect.scala 6:24]
  wire  fire_2 = idu_io_out_valid & issue_io_in_ready; // @[Connect.scala 7:27]
  wire  _T_5 = issue_io_in_ready & issue_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_26 = _T_5 ? 1'h0 : valid_2; // @[Connect.scala 8:23 Connect.scala 8:31 Connect.scala 6:24]
  wire  _GEN_27 = fire_2 | _GEN_26; // @[Connect.scala 9:17 Connect.scala 9:25]
  reg  issue_io_in_bits_r_0_valid; // @[Reg.scala 27:20]
  reg [31:0] issue_io_in_bits_r_0_pc; // @[Reg.scala 27:20]
  reg [31:0] issue_io_in_bits_r_0_inst; // @[Reg.scala 27:20]
  reg [1:0] issue_io_in_bits_r_0_src1; // @[Reg.scala 27:20]
  reg [1:0] issue_io_in_bits_r_0_src2; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_0_rs1; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_0_rs2; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_0_dest; // @[Reg.scala 27:20]
  reg [63:0] issue_io_in_bits_r_0_imm; // @[Reg.scala 27:20]
  reg [2:0] issue_io_in_bits_r_0_fu_type; // @[Reg.scala 27:20]
  reg [3:0] issue_io_in_bits_r_0_bru_op; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_0_alu_op; // @[Reg.scala 27:20]
  reg [3:0] issue_io_in_bits_r_0_lsu_op; // @[Reg.scala 27:20]
  reg [2:0] issue_io_in_bits_r_0_csr_op; // @[Reg.scala 27:20]
  reg [3:0] issue_io_in_bits_r_0_mdu_op; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_0_wen; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_0_rv64; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_0_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] issue_io_in_bits_r_0_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] issue_io_in_bits_r_0_bp_br_type; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_1_valid; // @[Reg.scala 27:20]
  reg [31:0] issue_io_in_bits_r_1_pc; // @[Reg.scala 27:20]
  reg [31:0] issue_io_in_bits_r_1_inst; // @[Reg.scala 27:20]
  reg [1:0] issue_io_in_bits_r_1_src1; // @[Reg.scala 27:20]
  reg [1:0] issue_io_in_bits_r_1_src2; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_1_rs1; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_1_rs2; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_1_dest; // @[Reg.scala 27:20]
  reg [63:0] issue_io_in_bits_r_1_imm; // @[Reg.scala 27:20]
  reg [2:0] issue_io_in_bits_r_1_fu_type; // @[Reg.scala 27:20]
  reg [3:0] issue_io_in_bits_r_1_bru_op; // @[Reg.scala 27:20]
  reg [4:0] issue_io_in_bits_r_1_alu_op; // @[Reg.scala 27:20]
  reg [3:0] issue_io_in_bits_r_1_lsu_op; // @[Reg.scala 27:20]
  reg [2:0] issue_io_in_bits_r_1_csr_op; // @[Reg.scala 27:20]
  reg [3:0] issue_io_in_bits_r_1_mdu_op; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_1_wen; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_1_rv64; // @[Reg.scala 27:20]
  reg  issue_io_in_bits_r_1_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] issue_io_in_bits_r_1_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] issue_io_in_bits_r_1_bp_br_type; // @[Reg.scala 27:20]
  reg  valid_3; // @[Connect.scala 6:24]
  wire  fire_3 = issue_io_out_valid & exu_io_in_ready; // @[Connect.scala 7:27]
  wire  _T_7 = exu_io_in_ready & exu_io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_69 = _T_7 ? 1'h0 : valid_3; // @[Connect.scala 8:23 Connect.scala 8:31 Connect.scala 6:24]
  wire  _GEN_70 = fire_3 | _GEN_69; // @[Connect.scala 9:17 Connect.scala 9:25]
  reg  exu_io_in_bits_r_0_valid; // @[Reg.scala 27:20]
  reg [31:0] exu_io_in_bits_r_0_pc; // @[Reg.scala 27:20]
  reg [31:0] exu_io_in_bits_r_0_inst; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_0_src1_value; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_0_src2_value; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_0_rs2_value; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_0_imm; // @[Reg.scala 27:20]
  reg [4:0] exu_io_in_bits_r_0_rs1; // @[Reg.scala 27:20]
  reg [4:0] exu_io_in_bits_r_0_dest; // @[Reg.scala 27:20]
  reg [2:0] exu_io_in_bits_r_0_fu_type; // @[Reg.scala 27:20]
  reg [3:0] exu_io_in_bits_r_0_bru_op; // @[Reg.scala 27:20]
  reg [4:0] exu_io_in_bits_r_0_alu_op; // @[Reg.scala 27:20]
  reg [3:0] exu_io_in_bits_r_0_lsu_op; // @[Reg.scala 27:20]
  reg [2:0] exu_io_in_bits_r_0_csr_op; // @[Reg.scala 27:20]
  reg [3:0] exu_io_in_bits_r_0_mdu_op; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_0_wen; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_0_rv64; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_0_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] exu_io_in_bits_r_0_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] exu_io_in_bits_r_0_bp_br_type; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_1_valid; // @[Reg.scala 27:20]
  reg [31:0] exu_io_in_bits_r_1_pc; // @[Reg.scala 27:20]
  reg [31:0] exu_io_in_bits_r_1_inst; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_1_src1_value; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_1_src2_value; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_1_rs2_value; // @[Reg.scala 27:20]
  reg [63:0] exu_io_in_bits_r_1_imm; // @[Reg.scala 27:20]
  reg [4:0] exu_io_in_bits_r_1_rs1; // @[Reg.scala 27:20]
  reg [4:0] exu_io_in_bits_r_1_dest; // @[Reg.scala 27:20]
  reg [2:0] exu_io_in_bits_r_1_fu_type; // @[Reg.scala 27:20]
  reg [3:0] exu_io_in_bits_r_1_bru_op; // @[Reg.scala 27:20]
  reg [4:0] exu_io_in_bits_r_1_alu_op; // @[Reg.scala 27:20]
  reg [3:0] exu_io_in_bits_r_1_lsu_op; // @[Reg.scala 27:20]
  reg [2:0] exu_io_in_bits_r_1_csr_op; // @[Reg.scala 27:20]
  reg [3:0] exu_io_in_bits_r_1_mdu_op; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_1_wen; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_1_rv64; // @[Reg.scala 27:20]
  reg  exu_io_in_bits_r_1_bp_br_taken; // @[Reg.scala 27:20]
  reg [31:0] exu_io_in_bits_r_1_bp_br_target; // @[Reg.scala 27:20]
  reg [1:0] exu_io_in_bits_r_1_bp_br_type; // @[Reg.scala 27:20]
  reg  valid_4; // @[Connect.scala 6:24]
  wire  fire_4 = exu_io_out_valid; // @[Connect.scala 7:27]
  wire  _T_8 = wbu_io__in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_112 = _T_8 ? 1'h0 : valid_4; // @[Connect.scala 8:23 Connect.scala 8:31 Connect.scala 6:24]
  wire  _GEN_113 = fire_4 | _GEN_112; // @[Connect.scala 9:17 Connect.scala 9:25]
  reg  wbu_io_in_bits_r_0_valid; // @[Reg.scala 27:20]
  reg [31:0] wbu_io_in_bits_r_0_pc; // @[Reg.scala 27:20]
  reg [63:0] wbu_io_in_bits_r_0_final_result; // @[Reg.scala 27:20]
  reg [4:0] wbu_io_in_bits_r_0_dest; // @[Reg.scala 27:20]
  reg  wbu_io_in_bits_r_0_wen; // @[Reg.scala 27:20]
  reg  wbu_io_in_bits_r_1_valid; // @[Reg.scala 27:20]
  reg [63:0] wbu_io_in_bits_r_1_final_result; // @[Reg.scala 27:20]
  reg [4:0] wbu_io_in_bits_r_1_dest; // @[Reg.scala 27:20]
  reg  wbu_io_in_bits_r_1_wen; // @[Reg.scala 27:20]
  IFU ifu ( // @[Core.scala 12:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_valid(ifu_io_imem_valid),
    .io_imem_addr(ifu_io_imem_addr),
    .io_imem_fence(ifu_io_imem_fence),
    .io_imem_fence_finish(ifu_io_imem_fence_finish),
    .io_imem_data_ok(ifu_io_imem_data_ok),
    .io_imem_inst(ifu_io_imem_inst),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_inst(ifu_io_out_bits_inst),
    .io_out_bits_uncache(ifu_io_out_bits_uncache),
    .io_out_bits_offset(ifu_io_out_bits_offset),
    .io_out_bits_bp_br_offset(ifu_io_out_bits_bp_br_offset),
    .io_out_bits_bp_br_taken(ifu_io_out_bits_bp_br_taken),
    .io_out_bits_bp_br_target(ifu_io_out_bits_bp_br_target),
    .io_out_bits_bp_br_type(ifu_io_out_bits_bp_br_type),
    .io_reflush_bus_is_reflush(ifu_io_reflush_bus_is_reflush),
    .io_reflush_bus_br_target(ifu_io_reflush_bus_br_target),
    .io_bpu_valid(ifu_io_bpu_valid),
    .io_bpu_pc(ifu_io_bpu_pc),
    .io_bpu_bp_ok(ifu_io_bpu_bp_ok),
    .io_bpu_bp_taken(ifu_io_bpu_bp_taken),
    .io_bpu_bp_target(ifu_io_bpu_bp_target),
    .io_bpu_bp_offset(ifu_io_bpu_bp_offset),
    .io_bpu_is_reflush(ifu_io_bpu_is_reflush),
    .io_bpu_bp_type(ifu_io_bpu_bp_type),
    .io_bpu_call_count(ifu_io_bpu_call_count),
    .io_bpu_ret_count(ifu_io_bpu_ret_count),
    .dcache_fence_finish_0(ifu_dcache_fence_finish_0),
    .fence_i(ifu_fence_i),
    .icache_fence_finish_0(ifu_icache_fence_finish_0)
  );
  IQueue iqueue ( // @[Core.scala 13:22]
    .clock(iqueue_clock),
    .reset(iqueue_reset),
    .io_in_ready(iqueue_io_in_ready),
    .io_in_valid(iqueue_io_in_valid),
    .io_in_bits_pc(iqueue_io_in_bits_pc),
    .io_in_bits_inst(iqueue_io_in_bits_inst),
    .io_in_bits_uncache(iqueue_io_in_bits_uncache),
    .io_in_bits_offset(iqueue_io_in_bits_offset),
    .io_in_bits_bp_br_offset(iqueue_io_in_bits_bp_br_offset),
    .io_in_bits_bp_br_taken(iqueue_io_in_bits_bp_br_taken),
    .io_in_bits_bp_br_target(iqueue_io_in_bits_bp_br_target),
    .io_in_bits_bp_br_type(iqueue_io_in_bits_bp_br_type),
    .io_out_ready(iqueue_io_out_ready),
    .io_out_valid(iqueue_io_out_valid),
    .io_out_bits_0_valid(iqueue_io_out_bits_0_valid),
    .io_out_bits_0_pc(iqueue_io_out_bits_0_pc),
    .io_out_bits_0_inst(iqueue_io_out_bits_0_inst),
    .io_out_bits_0_bp_br_taken(iqueue_io_out_bits_0_bp_br_taken),
    .io_out_bits_0_bp_br_target(iqueue_io_out_bits_0_bp_br_target),
    .io_out_bits_0_bp_br_type(iqueue_io_out_bits_0_bp_br_type),
    .io_out_bits_1_valid(iqueue_io_out_bits_1_valid),
    .io_out_bits_1_pc(iqueue_io_out_bits_1_pc),
    .io_out_bits_1_inst(iqueue_io_out_bits_1_inst),
    .io_out_bits_1_bp_br_taken(iqueue_io_out_bits_1_bp_br_taken),
    .io_out_bits_1_bp_br_target(iqueue_io_out_bits_1_bp_br_target),
    .io_out_bits_1_bp_br_type(iqueue_io_out_bits_1_bp_br_type),
    .frontend_reflush(iqueue_frontend_reflush)
  );
  IDU idu ( // @[Core.scala 14:19]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_in_ready(idu_io_in_ready),
    .io_in_valid(idu_io_in_valid),
    .io_in_bits_0_valid(idu_io_in_bits_0_valid),
    .io_in_bits_0_pc(idu_io_in_bits_0_pc),
    .io_in_bits_0_inst(idu_io_in_bits_0_inst),
    .io_in_bits_0_bp_br_taken(idu_io_in_bits_0_bp_br_taken),
    .io_in_bits_0_bp_br_target(idu_io_in_bits_0_bp_br_target),
    .io_in_bits_0_bp_br_type(idu_io_in_bits_0_bp_br_type),
    .io_in_bits_1_valid(idu_io_in_bits_1_valid),
    .io_in_bits_1_pc(idu_io_in_bits_1_pc),
    .io_in_bits_1_inst(idu_io_in_bits_1_inst),
    .io_in_bits_1_bp_br_taken(idu_io_in_bits_1_bp_br_taken),
    .io_in_bits_1_bp_br_target(idu_io_in_bits_1_bp_br_target),
    .io_in_bits_1_bp_br_type(idu_io_in_bits_1_bp_br_type),
    .io_out_ready(idu_io_out_ready),
    .io_out_valid(idu_io_out_valid),
    .io_out_bits_0_valid(idu_io_out_bits_0_valid),
    .io_out_bits_0_pc(idu_io_out_bits_0_pc),
    .io_out_bits_0_inst(idu_io_out_bits_0_inst),
    .io_out_bits_0_src1(idu_io_out_bits_0_src1),
    .io_out_bits_0_src2(idu_io_out_bits_0_src2),
    .io_out_bits_0_rs1(idu_io_out_bits_0_rs1),
    .io_out_bits_0_rs2(idu_io_out_bits_0_rs2),
    .io_out_bits_0_dest(idu_io_out_bits_0_dest),
    .io_out_bits_0_imm(idu_io_out_bits_0_imm),
    .io_out_bits_0_fu_type(idu_io_out_bits_0_fu_type),
    .io_out_bits_0_bru_op(idu_io_out_bits_0_bru_op),
    .io_out_bits_0_alu_op(idu_io_out_bits_0_alu_op),
    .io_out_bits_0_lsu_op(idu_io_out_bits_0_lsu_op),
    .io_out_bits_0_csr_op(idu_io_out_bits_0_csr_op),
    .io_out_bits_0_mdu_op(idu_io_out_bits_0_mdu_op),
    .io_out_bits_0_wen(idu_io_out_bits_0_wen),
    .io_out_bits_0_rv64(idu_io_out_bits_0_rv64),
    .io_out_bits_0_bp_br_taken(idu_io_out_bits_0_bp_br_taken),
    .io_out_bits_0_bp_br_target(idu_io_out_bits_0_bp_br_target),
    .io_out_bits_0_bp_br_type(idu_io_out_bits_0_bp_br_type),
    .io_out_bits_1_valid(idu_io_out_bits_1_valid),
    .io_out_bits_1_pc(idu_io_out_bits_1_pc),
    .io_out_bits_1_inst(idu_io_out_bits_1_inst),
    .io_out_bits_1_src1(idu_io_out_bits_1_src1),
    .io_out_bits_1_src2(idu_io_out_bits_1_src2),
    .io_out_bits_1_rs1(idu_io_out_bits_1_rs1),
    .io_out_bits_1_rs2(idu_io_out_bits_1_rs2),
    .io_out_bits_1_dest(idu_io_out_bits_1_dest),
    .io_out_bits_1_imm(idu_io_out_bits_1_imm),
    .io_out_bits_1_fu_type(idu_io_out_bits_1_fu_type),
    .io_out_bits_1_bru_op(idu_io_out_bits_1_bru_op),
    .io_out_bits_1_alu_op(idu_io_out_bits_1_alu_op),
    .io_out_bits_1_lsu_op(idu_io_out_bits_1_lsu_op),
    .io_out_bits_1_csr_op(idu_io_out_bits_1_csr_op),
    .io_out_bits_1_mdu_op(idu_io_out_bits_1_mdu_op),
    .io_out_bits_1_wen(idu_io_out_bits_1_wen),
    .io_out_bits_1_rv64(idu_io_out_bits_1_rv64),
    .io_out_bits_1_bp_br_taken(idu_io_out_bits_1_bp_br_taken),
    .io_out_bits_1_bp_br_target(idu_io_out_bits_1_bp_br_target),
    .io_out_bits_1_bp_br_type(idu_io_out_bits_1_bp_br_type),
    .frontend_reflush(idu_frontend_reflush)
  );
  Issue issue ( // @[Core.scala 15:21]
    .clock(issue_clock),
    .reset(issue_reset),
    .io_in_ready(issue_io_in_ready),
    .io_in_valid(issue_io_in_valid),
    .io_in_bits_0_valid(issue_io_in_bits_0_valid),
    .io_in_bits_0_pc(issue_io_in_bits_0_pc),
    .io_in_bits_0_inst(issue_io_in_bits_0_inst),
    .io_in_bits_0_src1(issue_io_in_bits_0_src1),
    .io_in_bits_0_src2(issue_io_in_bits_0_src2),
    .io_in_bits_0_rs1(issue_io_in_bits_0_rs1),
    .io_in_bits_0_rs2(issue_io_in_bits_0_rs2),
    .io_in_bits_0_dest(issue_io_in_bits_0_dest),
    .io_in_bits_0_imm(issue_io_in_bits_0_imm),
    .io_in_bits_0_fu_type(issue_io_in_bits_0_fu_type),
    .io_in_bits_0_bru_op(issue_io_in_bits_0_bru_op),
    .io_in_bits_0_alu_op(issue_io_in_bits_0_alu_op),
    .io_in_bits_0_lsu_op(issue_io_in_bits_0_lsu_op),
    .io_in_bits_0_csr_op(issue_io_in_bits_0_csr_op),
    .io_in_bits_0_mdu_op(issue_io_in_bits_0_mdu_op),
    .io_in_bits_0_wen(issue_io_in_bits_0_wen),
    .io_in_bits_0_rv64(issue_io_in_bits_0_rv64),
    .io_in_bits_0_bp_br_taken(issue_io_in_bits_0_bp_br_taken),
    .io_in_bits_0_bp_br_target(issue_io_in_bits_0_bp_br_target),
    .io_in_bits_0_bp_br_type(issue_io_in_bits_0_bp_br_type),
    .io_in_bits_1_valid(issue_io_in_bits_1_valid),
    .io_in_bits_1_pc(issue_io_in_bits_1_pc),
    .io_in_bits_1_inst(issue_io_in_bits_1_inst),
    .io_in_bits_1_src1(issue_io_in_bits_1_src1),
    .io_in_bits_1_src2(issue_io_in_bits_1_src2),
    .io_in_bits_1_rs1(issue_io_in_bits_1_rs1),
    .io_in_bits_1_rs2(issue_io_in_bits_1_rs2),
    .io_in_bits_1_dest(issue_io_in_bits_1_dest),
    .io_in_bits_1_imm(issue_io_in_bits_1_imm),
    .io_in_bits_1_fu_type(issue_io_in_bits_1_fu_type),
    .io_in_bits_1_bru_op(issue_io_in_bits_1_bru_op),
    .io_in_bits_1_alu_op(issue_io_in_bits_1_alu_op),
    .io_in_bits_1_lsu_op(issue_io_in_bits_1_lsu_op),
    .io_in_bits_1_csr_op(issue_io_in_bits_1_csr_op),
    .io_in_bits_1_mdu_op(issue_io_in_bits_1_mdu_op),
    .io_in_bits_1_wen(issue_io_in_bits_1_wen),
    .io_in_bits_1_rv64(issue_io_in_bits_1_rv64),
    .io_in_bits_1_bp_br_taken(issue_io_in_bits_1_bp_br_taken),
    .io_in_bits_1_bp_br_target(issue_io_in_bits_1_bp_br_target),
    .io_in_bits_1_bp_br_type(issue_io_in_bits_1_bp_br_type),
    .io_out_ready(issue_io_out_ready),
    .io_out_valid(issue_io_out_valid),
    .io_out_bits_0_valid(issue_io_out_bits_0_valid),
    .io_out_bits_0_pc(issue_io_out_bits_0_pc),
    .io_out_bits_0_inst(issue_io_out_bits_0_inst),
    .io_out_bits_0_src1_value(issue_io_out_bits_0_src1_value),
    .io_out_bits_0_src2_value(issue_io_out_bits_0_src2_value),
    .io_out_bits_0_rs2_value(issue_io_out_bits_0_rs2_value),
    .io_out_bits_0_imm(issue_io_out_bits_0_imm),
    .io_out_bits_0_rs1(issue_io_out_bits_0_rs1),
    .io_out_bits_0_dest(issue_io_out_bits_0_dest),
    .io_out_bits_0_fu_type(issue_io_out_bits_0_fu_type),
    .io_out_bits_0_bru_op(issue_io_out_bits_0_bru_op),
    .io_out_bits_0_alu_op(issue_io_out_bits_0_alu_op),
    .io_out_bits_0_lsu_op(issue_io_out_bits_0_lsu_op),
    .io_out_bits_0_csr_op(issue_io_out_bits_0_csr_op),
    .io_out_bits_0_mdu_op(issue_io_out_bits_0_mdu_op),
    .io_out_bits_0_wen(issue_io_out_bits_0_wen),
    .io_out_bits_0_rv64(issue_io_out_bits_0_rv64),
    .io_out_bits_0_bp_br_taken(issue_io_out_bits_0_bp_br_taken),
    .io_out_bits_0_bp_br_target(issue_io_out_bits_0_bp_br_target),
    .io_out_bits_0_bp_br_type(issue_io_out_bits_0_bp_br_type),
    .io_out_bits_1_valid(issue_io_out_bits_1_valid),
    .io_out_bits_1_pc(issue_io_out_bits_1_pc),
    .io_out_bits_1_inst(issue_io_out_bits_1_inst),
    .io_out_bits_1_src1_value(issue_io_out_bits_1_src1_value),
    .io_out_bits_1_src2_value(issue_io_out_bits_1_src2_value),
    .io_out_bits_1_rs2_value(issue_io_out_bits_1_rs2_value),
    .io_out_bits_1_imm(issue_io_out_bits_1_imm),
    .io_out_bits_1_rs1(issue_io_out_bits_1_rs1),
    .io_out_bits_1_dest(issue_io_out_bits_1_dest),
    .io_out_bits_1_fu_type(issue_io_out_bits_1_fu_type),
    .io_out_bits_1_bru_op(issue_io_out_bits_1_bru_op),
    .io_out_bits_1_alu_op(issue_io_out_bits_1_alu_op),
    .io_out_bits_1_lsu_op(issue_io_out_bits_1_lsu_op),
    .io_out_bits_1_csr_op(issue_io_out_bits_1_csr_op),
    .io_out_bits_1_mdu_op(issue_io_out_bits_1_mdu_op),
    .io_out_bits_1_wen(issue_io_out_bits_1_wen),
    .io_out_bits_1_rv64(issue_io_out_bits_1_rv64),
    .io_out_bits_1_bp_br_taken(issue_io_out_bits_1_bp_br_taken),
    .io_out_bits_1_bp_br_target(issue_io_out_bits_1_bp_br_target),
    .io_out_bits_1_bp_br_type(issue_io_out_bits_1_bp_br_type),
    .io_wb_bus_0_rf_wen(issue_io_wb_bus_0_rf_wen),
    .io_wb_bus_0_rf_waddr(issue_io_wb_bus_0_rf_waddr),
    .io_wb_bus_0_rf_wdata(issue_io_wb_bus_0_rf_wdata),
    .io_wb_bus_1_rf_wen(issue_io_wb_bus_1_rf_wen),
    .io_wb_bus_1_rf_waddr(issue_io_wb_bus_1_rf_waddr),
    .io_wb_bus_1_rf_wdata(issue_io_wb_bus_1_rf_wdata),
    .io_ex_fwd_0_blk_valid(issue_io_ex_fwd_0_blk_valid),
    .io_ex_fwd_0_fwd_valid(issue_io_ex_fwd_0_fwd_valid),
    .io_ex_fwd_0_rf_waddr(issue_io_ex_fwd_0_rf_waddr),
    .io_ex_fwd_0_rf_wdata(issue_io_ex_fwd_0_rf_wdata),
    .io_ex_fwd_1_blk_valid(issue_io_ex_fwd_1_blk_valid),
    .io_ex_fwd_1_fwd_valid(issue_io_ex_fwd_1_fwd_valid),
    .io_ex_fwd_1_rf_waddr(issue_io_ex_fwd_1_rf_waddr),
    .io_ex_fwd_1_rf_wdata(issue_io_ex_fwd_1_rf_wdata),
    .frontend_reflush(issue_frontend_reflush)
  );
  EXU exu ( // @[Core.scala 16:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_dmem_valid(exu_io_dmem_valid),
    .io_dmem_op(exu_io_dmem_op),
    .io_dmem_addr(exu_io_dmem_addr),
    .io_dmem_wstrb(exu_io_dmem_wstrb),
    .io_dmem_wdata(exu_io_dmem_wdata),
    .io_dmem_fence(exu_io_dmem_fence),
    .io_dmem_fence_finish(exu_io_dmem_fence_finish),
    .io_dmem_data_ok(exu_io_dmem_data_ok),
    .io_dmem_rdata(exu_io_dmem_rdata),
    .io_in_ready(exu_io_in_ready),
    .io_in_valid(exu_io_in_valid),
    .io_in_bits_0_valid(exu_io_in_bits_0_valid),
    .io_in_bits_0_pc(exu_io_in_bits_0_pc),
    .io_in_bits_0_inst(exu_io_in_bits_0_inst),
    .io_in_bits_0_src1_value(exu_io_in_bits_0_src1_value),
    .io_in_bits_0_src2_value(exu_io_in_bits_0_src2_value),
    .io_in_bits_0_rs2_value(exu_io_in_bits_0_rs2_value),
    .io_in_bits_0_imm(exu_io_in_bits_0_imm),
    .io_in_bits_0_rs1(exu_io_in_bits_0_rs1),
    .io_in_bits_0_dest(exu_io_in_bits_0_dest),
    .io_in_bits_0_fu_type(exu_io_in_bits_0_fu_type),
    .io_in_bits_0_bru_op(exu_io_in_bits_0_bru_op),
    .io_in_bits_0_alu_op(exu_io_in_bits_0_alu_op),
    .io_in_bits_0_lsu_op(exu_io_in_bits_0_lsu_op),
    .io_in_bits_0_csr_op(exu_io_in_bits_0_csr_op),
    .io_in_bits_0_mdu_op(exu_io_in_bits_0_mdu_op),
    .io_in_bits_0_wen(exu_io_in_bits_0_wen),
    .io_in_bits_0_rv64(exu_io_in_bits_0_rv64),
    .io_in_bits_0_bp_br_taken(exu_io_in_bits_0_bp_br_taken),
    .io_in_bits_0_bp_br_target(exu_io_in_bits_0_bp_br_target),
    .io_in_bits_0_bp_br_type(exu_io_in_bits_0_bp_br_type),
    .io_in_bits_1_valid(exu_io_in_bits_1_valid),
    .io_in_bits_1_pc(exu_io_in_bits_1_pc),
    .io_in_bits_1_inst(exu_io_in_bits_1_inst),
    .io_in_bits_1_src1_value(exu_io_in_bits_1_src1_value),
    .io_in_bits_1_src2_value(exu_io_in_bits_1_src2_value),
    .io_in_bits_1_rs2_value(exu_io_in_bits_1_rs2_value),
    .io_in_bits_1_imm(exu_io_in_bits_1_imm),
    .io_in_bits_1_rs1(exu_io_in_bits_1_rs1),
    .io_in_bits_1_dest(exu_io_in_bits_1_dest),
    .io_in_bits_1_fu_type(exu_io_in_bits_1_fu_type),
    .io_in_bits_1_bru_op(exu_io_in_bits_1_bru_op),
    .io_in_bits_1_alu_op(exu_io_in_bits_1_alu_op),
    .io_in_bits_1_lsu_op(exu_io_in_bits_1_lsu_op),
    .io_in_bits_1_csr_op(exu_io_in_bits_1_csr_op),
    .io_in_bits_1_mdu_op(exu_io_in_bits_1_mdu_op),
    .io_in_bits_1_wen(exu_io_in_bits_1_wen),
    .io_in_bits_1_rv64(exu_io_in_bits_1_rv64),
    .io_in_bits_1_bp_br_taken(exu_io_in_bits_1_bp_br_taken),
    .io_in_bits_1_bp_br_target(exu_io_in_bits_1_bp_br_target),
    .io_in_bits_1_bp_br_type(exu_io_in_bits_1_bp_br_type),
    .io_out_valid(exu_io_out_valid),
    .io_out_bits_0_valid(exu_io_out_bits_0_valid),
    .io_out_bits_0_pc(exu_io_out_bits_0_pc),
    .io_out_bits_0_final_result(exu_io_out_bits_0_final_result),
    .io_out_bits_0_dest(exu_io_out_bits_0_dest),
    .io_out_bits_0_wen(exu_io_out_bits_0_wen),
    .io_out_bits_1_valid(exu_io_out_bits_1_valid),
    .io_out_bits_1_final_result(exu_io_out_bits_1_final_result),
    .io_out_bits_1_dest(exu_io_out_bits_1_dest),
    .io_out_bits_1_wen(exu_io_out_bits_1_wen),
    .io_forward_0_blk_valid(exu_io_forward_0_blk_valid),
    .io_forward_0_fwd_valid(exu_io_forward_0_fwd_valid),
    .io_forward_0_rf_waddr(exu_io_forward_0_rf_waddr),
    .io_forward_0_rf_wdata(exu_io_forward_0_rf_wdata),
    .io_forward_1_blk_valid(exu_io_forward_1_blk_valid),
    .io_forward_1_fwd_valid(exu_io_forward_1_fwd_valid),
    .io_forward_1_rf_waddr(exu_io_forward_1_rf_waddr),
    .io_forward_1_rf_wdata(exu_io_forward_1_rf_wdata),
    .io_reflush_bus_is_reflush(exu_io_reflush_bus_is_reflush),
    .io_reflush_bus_br_target(exu_io_reflush_bus_br_target),
    .io_bpu_valid(exu_io_bpu_valid),
    .io_bpu_pc(exu_io_bpu_pc),
    .io_bpu_bp_taken(exu_io_bpu_bp_taken),
    .io_bpu_bp_target(exu_io_bpu_bp_target),
    .io_bpu_bp_type(exu_io_bpu_bp_type),
    .io_bpu_bp_wrong(exu_io_bpu_bp_wrong),
    .io_bpu_fence(exu_io_bpu_fence),
    .io_bpu_call_count(exu_io_bpu_call_count),
    .io_bpu_ret_count(exu_io_bpu_ret_count),
    .frontend_reflush_0(exu_frontend_reflush_0),
    .dcache_fence_finish(exu_dcache_fence_finish),
    .fence_0(exu_fence_0),
    .icache_fence_finish(exu_icache_fence_finish)
  );
  WBU wbu ( // @[Core.scala 17:19]
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_0_valid(wbu_io__in_bits_0_valid),
    .io__in_bits_0_pc(wbu_io__in_bits_0_pc),
    .io__in_bits_0_final_result(wbu_io__in_bits_0_final_result),
    .io__in_bits_0_dest(wbu_io__in_bits_0_dest),
    .io__in_bits_0_wen(wbu_io__in_bits_0_wen),
    .io__in_bits_1_valid(wbu_io__in_bits_1_valid),
    .io__in_bits_1_final_result(wbu_io__in_bits_1_final_result),
    .io__in_bits_1_dest(wbu_io__in_bits_1_dest),
    .io__in_bits_1_wen(wbu_io__in_bits_1_wen),
    .io__wb_bus_0_rf_wen(wbu_io__wb_bus_0_rf_wen),
    .io__wb_bus_0_rf_waddr(wbu_io__wb_bus_0_rf_waddr),
    .io__wb_bus_0_rf_wdata(wbu_io__wb_bus_0_rf_wdata),
    .io__wb_bus_1_rf_wen(wbu_io__wb_bus_1_rf_wen),
    .io__wb_bus_1_rf_waddr(wbu_io__wb_bus_1_rf_waddr),
    .io__wb_bus_1_rf_wdata(wbu_io__wb_bus_1_rf_wdata),
    .io__commit_0_pc(wbu_io__commit_0_pc),
    .io_commit_0_pc(wbu_io_commit_0_pc)
  );
  BPU bpu ( // @[Core.scala 18:19]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_ifu_valid(bpu_io_ifu_valid),
    .io_ifu_pc(bpu_io_ifu_pc),
    .io_ifu_bp_ok(bpu_io_ifu_bp_ok),
    .io_ifu_bp_taken(bpu_io_ifu_bp_taken),
    .io_ifu_bp_target(bpu_io_ifu_bp_target),
    .io_ifu_bp_offset(bpu_io_ifu_bp_offset),
    .io_ifu_is_reflush(bpu_io_ifu_is_reflush),
    .io_ifu_bp_type(bpu_io_ifu_bp_type),
    .io_ifu_call_count(bpu_io_ifu_call_count),
    .io_ifu_ret_count(bpu_io_ifu_ret_count),
    .io_exu_valid(bpu_io_exu_valid),
    .io_exu_pc(bpu_io_exu_pc),
    .io_exu_bp_taken(bpu_io_exu_bp_taken),
    .io_exu_bp_target(bpu_io_exu_bp_target),
    .io_exu_bp_type(bpu_io_exu_bp_type),
    .io_exu_bp_wrong(bpu_io_exu_bp_wrong),
    .io_exu_fence(bpu_io_exu_fence),
    .io_exu_call_count(bpu_io_exu_call_count),
    .io_exu_ret_count(bpu_io_exu_ret_count)
  );
  Cache_Soc icache ( // @[Core.scala 19:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_in_valid(icache_io_in_valid),
    .io_in_op(icache_io_in_op),
    .io_in_addr(icache_io_in_addr),
    .io_in_wstrb(icache_io_in_wstrb),
    .io_in_wdata(icache_io_in_wdata),
    .io_in_fence(icache_io_in_fence),
    .io_in_fence_finish(icache_io_in_fence_finish),
    .io_in_data_ok(icache_io_in_data_ok),
    .io_in_rdata(icache_io_in_rdata),
    .io_in_inst(icache_io_in_inst),
    .io_out_rd_req(icache_io_out_rd_req),
    .io_out_rd_size(icache_io_out_rd_size),
    .io_out_rd_addr(icache_io_out_rd_addr),
    .io_out_rd_rdy(icache_io_out_rd_rdy),
    .io_out_ret_valid(icache_io_out_ret_valid),
    .io_out_ret_data(icache_io_out_ret_data),
    .io_out_wr_req(icache_io_out_wr_req),
    .io_out_wr_size(icache_io_out_wr_size),
    .io_out_wr_addr(icache_io_out_wr_addr),
    .io_out_wr_wstrb(icache_io_out_wr_wstrb),
    .io_out_wr_data(icache_io_out_wr_data),
    .io_out_wr_rdy(icache_io_out_wr_rdy),
    .io_out_wr_ok(icache_io_out_wr_ok),
    .io_sram_0_en(icache_io_sram_0_en),
    .io_sram_0_wen(icache_io_sram_0_wen),
    .io_sram_0_addr(icache_io_sram_0_addr),
    .io_sram_0_wdata(icache_io_sram_0_wdata),
    .io_sram_0_rdata(icache_io_sram_0_rdata),
    .io_sram_1_en(icache_io_sram_1_en),
    .io_sram_1_wen(icache_io_sram_1_wen),
    .io_sram_1_addr(icache_io_sram_1_addr),
    .io_sram_1_wdata(icache_io_sram_1_wdata),
    .io_sram_1_rdata(icache_io_sram_1_rdata),
    .io_sram_2_en(icache_io_sram_2_en),
    .io_sram_2_wen(icache_io_sram_2_wen),
    .io_sram_2_addr(icache_io_sram_2_addr),
    .io_sram_2_wdata(icache_io_sram_2_wdata),
    .io_sram_2_rdata(icache_io_sram_2_rdata),
    .io_sram_3_en(icache_io_sram_3_en),
    .io_sram_3_wen(icache_io_sram_3_wen),
    .io_sram_3_addr(icache_io_sram_3_addr),
    .io_sram_3_wdata(icache_io_sram_3_wdata),
    .io_sram_3_rdata(icache_io_sram_3_rdata)
  );
  Cache_Soc dcache ( // @[Core.scala 20:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_in_valid(dcache_io_in_valid),
    .io_in_op(dcache_io_in_op),
    .io_in_addr(dcache_io_in_addr),
    .io_in_wstrb(dcache_io_in_wstrb),
    .io_in_wdata(dcache_io_in_wdata),
    .io_in_fence(dcache_io_in_fence),
    .io_in_fence_finish(dcache_io_in_fence_finish),
    .io_in_data_ok(dcache_io_in_data_ok),
    .io_in_rdata(dcache_io_in_rdata),
    .io_in_inst(dcache_io_in_inst),
    .io_out_rd_req(dcache_io_out_rd_req),
    .io_out_rd_size(dcache_io_out_rd_size),
    .io_out_rd_addr(dcache_io_out_rd_addr),
    .io_out_rd_rdy(dcache_io_out_rd_rdy),
    .io_out_ret_valid(dcache_io_out_ret_valid),
    .io_out_ret_data(dcache_io_out_ret_data),
    .io_out_wr_req(dcache_io_out_wr_req),
    .io_out_wr_size(dcache_io_out_wr_size),
    .io_out_wr_addr(dcache_io_out_wr_addr),
    .io_out_wr_wstrb(dcache_io_out_wr_wstrb),
    .io_out_wr_data(dcache_io_out_wr_data),
    .io_out_wr_rdy(dcache_io_out_wr_rdy),
    .io_out_wr_ok(dcache_io_out_wr_ok),
    .io_sram_0_en(dcache_io_sram_0_en),
    .io_sram_0_wen(dcache_io_sram_0_wen),
    .io_sram_0_addr(dcache_io_sram_0_addr),
    .io_sram_0_wdata(dcache_io_sram_0_wdata),
    .io_sram_0_rdata(dcache_io_sram_0_rdata),
    .io_sram_1_en(dcache_io_sram_1_en),
    .io_sram_1_wen(dcache_io_sram_1_wen),
    .io_sram_1_addr(dcache_io_sram_1_addr),
    .io_sram_1_wdata(dcache_io_sram_1_wdata),
    .io_sram_1_rdata(dcache_io_sram_1_rdata),
    .io_sram_2_en(dcache_io_sram_2_en),
    .io_sram_2_wen(dcache_io_sram_2_wen),
    .io_sram_2_addr(dcache_io_sram_2_addr),
    .io_sram_2_wdata(dcache_io_sram_2_wdata),
    .io_sram_2_rdata(dcache_io_sram_2_rdata),
    .io_sram_3_en(dcache_io_sram_3_en),
    .io_sram_3_wen(dcache_io_sram_3_wen),
    .io_sram_3_addr(dcache_io_sram_3_addr),
    .io_sram_3_wdata(dcache_io_sram_3_wdata),
    .io_sram_3_rdata(dcache_io_sram_3_rdata)
  );
  assign io_icache_bridge_rd_req = icache_io_out_rd_req; // @[Core.scala 26:17]
  assign io_icache_bridge_rd_size = icache_io_out_rd_size; // @[Core.scala 26:17]
  assign io_icache_bridge_rd_addr = icache_io_out_rd_addr; // @[Core.scala 26:17]
  assign io_dcache_bridge_rd_req = dcache_io_out_rd_req; // @[Core.scala 39:17]
  assign io_dcache_bridge_rd_size = dcache_io_out_rd_size; // @[Core.scala 39:17]
  assign io_dcache_bridge_rd_addr = dcache_io_out_rd_addr; // @[Core.scala 39:17]
  assign io_dcache_bridge_wr_req = dcache_io_out_wr_req; // @[Core.scala 39:17]
  assign io_dcache_bridge_wr_size = dcache_io_out_wr_size; // @[Core.scala 39:17]
  assign io_dcache_bridge_wr_addr = dcache_io_out_wr_addr; // @[Core.scala 39:17]
  assign io_dcache_bridge_wr_wstrb = dcache_io_out_wr_wstrb; // @[Core.scala 39:17]
  assign io_dcache_bridge_wr_data = dcache_io_out_wr_data; // @[Core.scala 39:17]
  assign io_sram_0_en = icache_io_sram_0_en; // @[Core.scala 21:11]
  assign io_sram_0_wen = icache_io_sram_0_wen; // @[Core.scala 21:11]
  assign io_sram_0_addr = icache_io_sram_0_addr; // @[Core.scala 21:11]
  assign io_sram_0_wdata = icache_io_sram_0_wdata; // @[Core.scala 21:11]
  assign io_sram_1_en = icache_io_sram_1_en; // @[Core.scala 21:11]
  assign io_sram_1_wen = icache_io_sram_1_wen; // @[Core.scala 21:11]
  assign io_sram_1_addr = icache_io_sram_1_addr; // @[Core.scala 21:11]
  assign io_sram_1_wdata = icache_io_sram_1_wdata; // @[Core.scala 21:11]
  assign io_sram_2_en = icache_io_sram_2_en; // @[Core.scala 21:11]
  assign io_sram_2_wen = icache_io_sram_2_wen; // @[Core.scala 21:11]
  assign io_sram_2_addr = icache_io_sram_2_addr; // @[Core.scala 21:11]
  assign io_sram_2_wdata = icache_io_sram_2_wdata; // @[Core.scala 21:11]
  assign io_sram_3_en = icache_io_sram_3_en; // @[Core.scala 21:11]
  assign io_sram_3_wen = icache_io_sram_3_wen; // @[Core.scala 21:11]
  assign io_sram_3_addr = icache_io_sram_3_addr; // @[Core.scala 21:11]
  assign io_sram_3_wdata = icache_io_sram_3_wdata; // @[Core.scala 21:11]
  assign io_sram_4_en = dcache_io_sram_0_en; // @[Core.scala 21:11]
  assign io_sram_4_wen = dcache_io_sram_0_wen; // @[Core.scala 21:11]
  assign io_sram_4_addr = dcache_io_sram_0_addr; // @[Core.scala 21:11]
  assign io_sram_4_wdata = dcache_io_sram_0_wdata; // @[Core.scala 21:11]
  assign io_sram_5_en = dcache_io_sram_1_en; // @[Core.scala 21:11]
  assign io_sram_5_wen = dcache_io_sram_1_wen; // @[Core.scala 21:11]
  assign io_sram_5_addr = dcache_io_sram_1_addr; // @[Core.scala 21:11]
  assign io_sram_5_wdata = dcache_io_sram_1_wdata; // @[Core.scala 21:11]
  assign io_sram_6_en = dcache_io_sram_2_en; // @[Core.scala 21:11]
  assign io_sram_6_wen = dcache_io_sram_2_wen; // @[Core.scala 21:11]
  assign io_sram_6_addr = dcache_io_sram_2_addr; // @[Core.scala 21:11]
  assign io_sram_6_wdata = dcache_io_sram_2_wdata; // @[Core.scala 21:11]
  assign io_sram_7_en = dcache_io_sram_3_en; // @[Core.scala 21:11]
  assign io_sram_7_wen = dcache_io_sram_3_wen; // @[Core.scala 21:11]
  assign io_sram_7_addr = dcache_io_sram_3_addr; // @[Core.scala 21:11]
  assign io_sram_7_wdata = dcache_io_sram_3_wdata; // @[Core.scala 21:11]
  assign io_commit_0_pc = wbu_io_commit_0_pc;
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_fence_finish = icache_io_in_fence_finish; // @[Core.scala 27:15]
  assign ifu_io_imem_data_ok = icache_io_in_data_ok; // @[Core.scala 27:15]
  assign ifu_io_imem_inst = icache_io_in_inst; // @[Core.scala 27:15]
  assign ifu_io_out_ready = iqueue_io_in_ready; // @[Connect.scala 12:16]
  assign ifu_io_reflush_bus_is_reflush = exu_io_reflush_bus_is_reflush; // @[Core.scala 28:22]
  assign ifu_io_reflush_bus_br_target = exu_io_reflush_bus_br_target; // @[Core.scala 28:22]
  assign ifu_io_bpu_bp_ok = bpu_io_ifu_bp_ok; // @[Core.scala 29:14]
  assign ifu_io_bpu_bp_taken = bpu_io_ifu_bp_taken; // @[Core.scala 29:14]
  assign ifu_io_bpu_bp_target = bpu_io_ifu_bp_target; // @[Core.scala 29:14]
  assign ifu_io_bpu_bp_offset = bpu_io_ifu_bp_offset; // @[Core.scala 29:14]
  assign ifu_io_bpu_bp_type = bpu_io_ifu_bp_type; // @[Core.scala 29:14]
  assign ifu_dcache_fence_finish_0 = exu_dcache_fence_finish;
  assign ifu_fence_i = exu_fence_0;
  assign iqueue_clock = clock;
  assign iqueue_reset = reset;
  assign iqueue_io_in_valid = valid; // @[Connect.scala 14:17]
  assign iqueue_io_in_bits_pc = iqueue_io_in_bits_r_pc; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_inst = iqueue_io_in_bits_r_inst; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_uncache = iqueue_io_in_bits_r_uncache; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_offset = iqueue_io_in_bits_r_offset; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_bp_br_offset = iqueue_io_in_bits_r_bp_br_offset; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_bp_br_taken = iqueue_io_in_bits_r_bp_br_taken; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_bp_br_target = iqueue_io_in_bits_r_bp_br_target; // @[Connect.scala 13:16]
  assign iqueue_io_in_bits_bp_br_type = iqueue_io_in_bits_r_bp_br_type; // @[Connect.scala 13:16]
  assign iqueue_io_out_ready = idu_io_in_ready; // @[Connect.scala 12:16]
  assign iqueue_frontend_reflush = exu_frontend_reflush_0;
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_in_valid = valid_1; // @[Connect.scala 14:17]
  assign idu_io_in_bits_0_valid = idu_io_in_bits_r_0_valid; // @[Connect.scala 13:16]
  assign idu_io_in_bits_0_pc = idu_io_in_bits_r_0_pc; // @[Connect.scala 13:16]
  assign idu_io_in_bits_0_inst = idu_io_in_bits_r_0_inst; // @[Connect.scala 13:16]
  assign idu_io_in_bits_0_bp_br_taken = idu_io_in_bits_r_0_bp_br_taken; // @[Connect.scala 13:16]
  assign idu_io_in_bits_0_bp_br_target = idu_io_in_bits_r_0_bp_br_target; // @[Connect.scala 13:16]
  assign idu_io_in_bits_0_bp_br_type = idu_io_in_bits_r_0_bp_br_type; // @[Connect.scala 13:16]
  assign idu_io_in_bits_1_valid = idu_io_in_bits_r_1_valid; // @[Connect.scala 13:16]
  assign idu_io_in_bits_1_pc = idu_io_in_bits_r_1_pc; // @[Connect.scala 13:16]
  assign idu_io_in_bits_1_inst = idu_io_in_bits_r_1_inst; // @[Connect.scala 13:16]
  assign idu_io_in_bits_1_bp_br_taken = idu_io_in_bits_r_1_bp_br_taken; // @[Connect.scala 13:16]
  assign idu_io_in_bits_1_bp_br_target = idu_io_in_bits_r_1_bp_br_target; // @[Connect.scala 13:16]
  assign idu_io_in_bits_1_bp_br_type = idu_io_in_bits_r_1_bp_br_type; // @[Connect.scala 13:16]
  assign idu_io_out_ready = issue_io_in_ready; // @[Connect.scala 12:16]
  assign idu_frontend_reflush = exu_frontend_reflush_0;
  assign issue_clock = clock;
  assign issue_reset = reset;
  assign issue_io_in_valid = valid_2; // @[Connect.scala 14:17]
  assign issue_io_in_bits_0_valid = issue_io_in_bits_r_0_valid; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_pc = issue_io_in_bits_r_0_pc; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_inst = issue_io_in_bits_r_0_inst; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_src1 = issue_io_in_bits_r_0_src1; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_src2 = issue_io_in_bits_r_0_src2; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_rs1 = issue_io_in_bits_r_0_rs1; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_rs2 = issue_io_in_bits_r_0_rs2; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_dest = issue_io_in_bits_r_0_dest; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_imm = issue_io_in_bits_r_0_imm; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_fu_type = issue_io_in_bits_r_0_fu_type; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_bru_op = issue_io_in_bits_r_0_bru_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_alu_op = issue_io_in_bits_r_0_alu_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_lsu_op = issue_io_in_bits_r_0_lsu_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_csr_op = issue_io_in_bits_r_0_csr_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_mdu_op = issue_io_in_bits_r_0_mdu_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_wen = issue_io_in_bits_r_0_wen; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_rv64 = issue_io_in_bits_r_0_rv64; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_bp_br_taken = issue_io_in_bits_r_0_bp_br_taken; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_bp_br_target = issue_io_in_bits_r_0_bp_br_target; // @[Connect.scala 13:16]
  assign issue_io_in_bits_0_bp_br_type = issue_io_in_bits_r_0_bp_br_type; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_valid = issue_io_in_bits_r_1_valid; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_pc = issue_io_in_bits_r_1_pc; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_inst = issue_io_in_bits_r_1_inst; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_src1 = issue_io_in_bits_r_1_src1; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_src2 = issue_io_in_bits_r_1_src2; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_rs1 = issue_io_in_bits_r_1_rs1; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_rs2 = issue_io_in_bits_r_1_rs2; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_dest = issue_io_in_bits_r_1_dest; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_imm = issue_io_in_bits_r_1_imm; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_fu_type = issue_io_in_bits_r_1_fu_type; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_bru_op = issue_io_in_bits_r_1_bru_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_alu_op = issue_io_in_bits_r_1_alu_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_lsu_op = issue_io_in_bits_r_1_lsu_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_csr_op = issue_io_in_bits_r_1_csr_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_mdu_op = issue_io_in_bits_r_1_mdu_op; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_wen = issue_io_in_bits_r_1_wen; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_rv64 = issue_io_in_bits_r_1_rv64; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_bp_br_taken = issue_io_in_bits_r_1_bp_br_taken; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_bp_br_target = issue_io_in_bits_r_1_bp_br_target; // @[Connect.scala 13:16]
  assign issue_io_in_bits_1_bp_br_type = issue_io_in_bits_r_1_bp_br_type; // @[Connect.scala 13:16]
  assign issue_io_out_ready = exu_io_in_ready; // @[Connect.scala 12:16]
  assign issue_io_wb_bus_0_rf_wen = wbu_io__wb_bus_0_rf_wen; // @[Core.scala 34:19]
  assign issue_io_wb_bus_0_rf_waddr = wbu_io__wb_bus_0_rf_waddr; // @[Core.scala 34:19]
  assign issue_io_wb_bus_0_rf_wdata = wbu_io__wb_bus_0_rf_wdata; // @[Core.scala 34:19]
  assign issue_io_wb_bus_1_rf_wen = wbu_io__wb_bus_1_rf_wen; // @[Core.scala 34:19]
  assign issue_io_wb_bus_1_rf_waddr = wbu_io__wb_bus_1_rf_waddr; // @[Core.scala 34:19]
  assign issue_io_wb_bus_1_rf_wdata = wbu_io__wb_bus_1_rf_wdata; // @[Core.scala 34:19]
  assign issue_io_ex_fwd_0_blk_valid = exu_io_forward_0_blk_valid; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_0_fwd_valid = exu_io_forward_0_fwd_valid; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_0_rf_waddr = exu_io_forward_0_rf_waddr; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_0_rf_wdata = exu_io_forward_0_rf_wdata; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_1_blk_valid = exu_io_forward_1_blk_valid; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_1_fwd_valid = exu_io_forward_1_fwd_valid; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_1_rf_waddr = exu_io_forward_1_rf_waddr; // @[Core.scala 35:19]
  assign issue_io_ex_fwd_1_rf_wdata = exu_io_forward_1_rf_wdata; // @[Core.scala 35:19]
  assign issue_frontend_reflush = exu_frontend_reflush_0;
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_dmem_fence_finish = dcache_io_in_fence_finish; // @[Core.scala 40:15]
  assign exu_io_dmem_data_ok = dcache_io_in_data_ok; // @[Core.scala 40:15]
  assign exu_io_dmem_rdata = dcache_io_in_rdata; // @[Core.scala 40:15]
  assign exu_io_in_valid = valid_3; // @[Connect.scala 14:17]
  assign exu_io_in_bits_0_valid = exu_io_in_bits_r_0_valid; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_pc = exu_io_in_bits_r_0_pc; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_inst = exu_io_in_bits_r_0_inst; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_src1_value = exu_io_in_bits_r_0_src1_value; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_src2_value = exu_io_in_bits_r_0_src2_value; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_rs2_value = exu_io_in_bits_r_0_rs2_value; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_imm = exu_io_in_bits_r_0_imm; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_rs1 = exu_io_in_bits_r_0_rs1; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_dest = exu_io_in_bits_r_0_dest; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_fu_type = exu_io_in_bits_r_0_fu_type; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_bru_op = exu_io_in_bits_r_0_bru_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_alu_op = exu_io_in_bits_r_0_alu_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_lsu_op = exu_io_in_bits_r_0_lsu_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_csr_op = exu_io_in_bits_r_0_csr_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_mdu_op = exu_io_in_bits_r_0_mdu_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_wen = exu_io_in_bits_r_0_wen; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_rv64 = exu_io_in_bits_r_0_rv64; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_bp_br_taken = exu_io_in_bits_r_0_bp_br_taken; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_bp_br_target = exu_io_in_bits_r_0_bp_br_target; // @[Connect.scala 13:16]
  assign exu_io_in_bits_0_bp_br_type = exu_io_in_bits_r_0_bp_br_type; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_valid = exu_io_in_bits_r_1_valid; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_pc = exu_io_in_bits_r_1_pc; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_inst = exu_io_in_bits_r_1_inst; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_src1_value = exu_io_in_bits_r_1_src1_value; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_src2_value = exu_io_in_bits_r_1_src2_value; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_rs2_value = exu_io_in_bits_r_1_rs2_value; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_imm = exu_io_in_bits_r_1_imm; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_rs1 = exu_io_in_bits_r_1_rs1; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_dest = exu_io_in_bits_r_1_dest; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_fu_type = exu_io_in_bits_r_1_fu_type; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_bru_op = exu_io_in_bits_r_1_bru_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_alu_op = exu_io_in_bits_r_1_alu_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_lsu_op = exu_io_in_bits_r_1_lsu_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_csr_op = exu_io_in_bits_r_1_csr_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_mdu_op = exu_io_in_bits_r_1_mdu_op; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_wen = exu_io_in_bits_r_1_wen; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_rv64 = exu_io_in_bits_r_1_rv64; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_bp_br_taken = exu_io_in_bits_r_1_bp_br_taken; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_bp_br_target = exu_io_in_bits_r_1_bp_br_target; // @[Connect.scala 13:16]
  assign exu_io_in_bits_1_bp_br_type = exu_io_in_bits_r_1_bp_br_type; // @[Connect.scala 13:16]
  assign exu_icache_fence_finish = ifu_icache_fence_finish_0;
  assign wbu_io__in_valid = valid_4; // @[Connect.scala 14:17]
  assign wbu_io__in_bits_0_valid = wbu_io_in_bits_r_0_valid; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_0_pc = wbu_io_in_bits_r_0_pc; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_0_final_result = wbu_io_in_bits_r_0_final_result; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_0_dest = wbu_io_in_bits_r_0_dest; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_0_wen = wbu_io_in_bits_r_0_wen; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_1_valid = wbu_io_in_bits_r_1_valid; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_1_final_result = wbu_io_in_bits_r_1_final_result; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_1_dest = wbu_io_in_bits_r_1_dest; // @[Connect.scala 13:16]
  assign wbu_io__in_bits_1_wen = wbu_io_in_bits_r_1_wen; // @[Connect.scala 13:16]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_ifu_valid = ifu_io_bpu_valid; // @[Core.scala 29:14]
  assign bpu_io_ifu_pc = ifu_io_bpu_pc; // @[Core.scala 29:14]
  assign bpu_io_ifu_is_reflush = ifu_io_bpu_is_reflush; // @[Core.scala 29:14]
  assign bpu_io_ifu_call_count = ifu_io_bpu_call_count; // @[Core.scala 29:14]
  assign bpu_io_ifu_ret_count = ifu_io_bpu_ret_count; // @[Core.scala 29:14]
  assign bpu_io_exu_valid = exu_io_bpu_valid; // @[Core.scala 41:14]
  assign bpu_io_exu_pc = exu_io_bpu_pc; // @[Core.scala 41:14]
  assign bpu_io_exu_bp_taken = exu_io_bpu_bp_taken; // @[Core.scala 41:14]
  assign bpu_io_exu_bp_target = exu_io_bpu_bp_target; // @[Core.scala 41:14]
  assign bpu_io_exu_bp_type = exu_io_bpu_bp_type; // @[Core.scala 41:14]
  assign bpu_io_exu_bp_wrong = exu_io_bpu_bp_wrong; // @[Core.scala 41:14]
  assign bpu_io_exu_fence = exu_io_bpu_fence; // @[Core.scala 41:14]
  assign bpu_io_exu_call_count = exu_io_bpu_call_count; // @[Core.scala 41:14]
  assign bpu_io_exu_ret_count = exu_io_bpu_ret_count; // @[Core.scala 41:14]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_in_valid = ifu_io_imem_valid; // @[Core.scala 27:15]
  assign icache_io_in_op = 1'h0; // @[Core.scala 27:15]
  assign icache_io_in_addr = ifu_io_imem_addr; // @[Core.scala 27:15]
  assign icache_io_in_wstrb = 8'h0; // @[Core.scala 27:15]
  assign icache_io_in_wdata = 64'h0; // @[Core.scala 27:15]
  assign icache_io_in_fence = ifu_io_imem_fence; // @[Core.scala 27:15]
  assign icache_io_out_rd_rdy = io_icache_bridge_rd_rdy; // @[Core.scala 26:17]
  assign icache_io_out_ret_valid = io_icache_bridge_ret_valid; // @[Core.scala 26:17]
  assign icache_io_out_ret_data = io_icache_bridge_ret_data; // @[Core.scala 26:17]
  assign icache_io_out_wr_rdy = 1'h1; // @[Core.scala 26:17]
  assign icache_io_out_wr_ok = 1'h1; // @[Core.scala 26:17]
  assign icache_io_sram_0_rdata = io_sram_0_rdata; // @[Core.scala 21:11]
  assign icache_io_sram_1_rdata = io_sram_1_rdata; // @[Core.scala 21:11]
  assign icache_io_sram_2_rdata = io_sram_2_rdata; // @[Core.scala 21:11]
  assign icache_io_sram_3_rdata = io_sram_3_rdata; // @[Core.scala 21:11]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_in_valid = exu_io_dmem_valid; // @[Core.scala 40:15]
  assign dcache_io_in_op = exu_io_dmem_op; // @[Core.scala 40:15]
  assign dcache_io_in_addr = exu_io_dmem_addr; // @[Core.scala 40:15]
  assign dcache_io_in_wstrb = exu_io_dmem_wstrb; // @[Core.scala 40:15]
  assign dcache_io_in_wdata = exu_io_dmem_wdata; // @[Core.scala 40:15]
  assign dcache_io_in_fence = exu_io_dmem_fence; // @[Core.scala 40:15]
  assign dcache_io_out_rd_rdy = io_dcache_bridge_rd_rdy; // @[Core.scala 39:17]
  assign dcache_io_out_ret_valid = io_dcache_bridge_ret_valid; // @[Core.scala 39:17]
  assign dcache_io_out_ret_data = io_dcache_bridge_ret_data; // @[Core.scala 39:17]
  assign dcache_io_out_wr_rdy = io_dcache_bridge_wr_rdy; // @[Core.scala 39:17]
  assign dcache_io_out_wr_ok = io_dcache_bridge_wr_ok; // @[Core.scala 39:17]
  assign dcache_io_sram_0_rdata = io_sram_4_rdata; // @[Core.scala 21:11]
  assign dcache_io_sram_1_rdata = io_sram_5_rdata; // @[Core.scala 21:11]
  assign dcache_io_sram_2_rdata = io_sram_6_rdata; // @[Core.scala 21:11]
  assign dcache_io_sram_3_rdata = io_sram_7_rdata; // @[Core.scala 21:11]
  always @(posedge clock) begin
    if (reset) begin // @[Connect.scala 6:24]
      valid <= 1'h0; // @[Connect.scala 6:24]
    end else if (frontend_reflush_0) begin // @[Connect.scala 10:23]
      valid <= 1'h0; // @[Connect.scala 10:30]
    end else begin
      valid <= _GEN_1;
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_pc <= ifu_io_out_bits_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_inst <= 128'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_inst <= ifu_io_out_bits_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_uncache <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_uncache <= ifu_io_out_bits_uncache; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_offset <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_offset <= ifu_io_out_bits_offset; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_bp_br_offset <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_bp_br_offset <= ifu_io_out_bits_bp_br_offset; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_bp_br_taken <= ifu_io_out_bits_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_bp_br_target <= ifu_io_out_bits_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      iqueue_io_in_bits_r_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire) begin // @[Reg.scala 28:19]
      iqueue_io_in_bits_r_bp_br_type <= ifu_io_out_bits_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Connect.scala 6:24]
      valid_1 <= 1'h0; // @[Connect.scala 6:24]
    end else if (frontend_reflush_0) begin // @[Connect.scala 10:23]
      valid_1 <= 1'h0; // @[Connect.scala 10:30]
    end else begin
      valid_1 <= _GEN_12;
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_0_valid <= iqueue_io_out_bits_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_0_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_0_pc <= iqueue_io_out_bits_0_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_0_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_0_inst <= iqueue_io_out_bits_0_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_0_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_0_bp_br_taken <= iqueue_io_out_bits_0_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_0_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_0_bp_br_target <= iqueue_io_out_bits_0_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_0_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_0_bp_br_type <= iqueue_io_out_bits_0_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_1_valid <= iqueue_io_out_bits_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_1_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_1_pc <= iqueue_io_out_bits_1_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_1_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_1_inst <= iqueue_io_out_bits_1_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_1_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_1_bp_br_taken <= iqueue_io_out_bits_1_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_1_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_1_bp_br_target <= iqueue_io_out_bits_1_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      idu_io_in_bits_r_1_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_1) begin // @[Reg.scala 28:19]
      idu_io_in_bits_r_1_bp_br_type <= iqueue_io_out_bits_1_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Connect.scala 6:24]
      valid_2 <= 1'h0; // @[Connect.scala 6:24]
    end else if (frontend_reflush_0) begin // @[Connect.scala 10:23]
      valid_2 <= 1'h0; // @[Connect.scala 10:30]
    end else begin
      valid_2 <= _GEN_27;
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_valid <= idu_io_out_bits_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_pc <= idu_io_out_bits_0_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_inst <= idu_io_out_bits_0_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_src1 <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_src1 <= idu_io_out_bits_0_src1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_src2 <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_src2 <= idu_io_out_bits_0_src2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_rs1 <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_rs1 <= idu_io_out_bits_0_rs1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_rs2 <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_rs2 <= idu_io_out_bits_0_rs2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_dest <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_dest <= idu_io_out_bits_0_dest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_imm <= idu_io_out_bits_0_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_fu_type <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_fu_type <= idu_io_out_bits_0_fu_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_bru_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_bru_op <= idu_io_out_bits_0_bru_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_alu_op <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_alu_op <= idu_io_out_bits_0_alu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_lsu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_lsu_op <= idu_io_out_bits_0_lsu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_csr_op <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_csr_op <= idu_io_out_bits_0_csr_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_mdu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_mdu_op <= idu_io_out_bits_0_mdu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_wen <= idu_io_out_bits_0_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_rv64 <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_rv64 <= idu_io_out_bits_0_rv64; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_bp_br_taken <= idu_io_out_bits_0_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_bp_br_target <= idu_io_out_bits_0_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_0_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_0_bp_br_type <= idu_io_out_bits_0_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_valid <= idu_io_out_bits_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_pc <= idu_io_out_bits_1_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_inst <= idu_io_out_bits_1_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_src1 <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_src1 <= idu_io_out_bits_1_src1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_src2 <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_src2 <= idu_io_out_bits_1_src2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_rs1 <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_rs1 <= idu_io_out_bits_1_rs1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_rs2 <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_rs2 <= idu_io_out_bits_1_rs2; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_dest <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_dest <= idu_io_out_bits_1_dest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_imm <= idu_io_out_bits_1_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_fu_type <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_fu_type <= idu_io_out_bits_1_fu_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_bru_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_bru_op <= idu_io_out_bits_1_bru_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_alu_op <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_alu_op <= idu_io_out_bits_1_alu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_lsu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_lsu_op <= idu_io_out_bits_1_lsu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_csr_op <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_csr_op <= idu_io_out_bits_1_csr_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_mdu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_mdu_op <= idu_io_out_bits_1_mdu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_wen <= idu_io_out_bits_1_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_rv64 <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_rv64 <= idu_io_out_bits_1_rv64; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_bp_br_taken <= idu_io_out_bits_1_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_bp_br_target <= idu_io_out_bits_1_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      issue_io_in_bits_r_1_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_2) begin // @[Reg.scala 28:19]
      issue_io_in_bits_r_1_bp_br_type <= idu_io_out_bits_1_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Connect.scala 6:24]
      valid_3 <= 1'h0; // @[Connect.scala 6:24]
    end else if (frontend_reflush_0) begin // @[Connect.scala 10:23]
      valid_3 <= 1'h0; // @[Connect.scala 10:30]
    end else begin
      valid_3 <= _GEN_70;
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_valid <= issue_io_out_bits_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_pc <= issue_io_out_bits_0_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_inst <= issue_io_out_bits_0_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_src1_value <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_src1_value <= issue_io_out_bits_0_src1_value; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_src2_value <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_src2_value <= issue_io_out_bits_0_src2_value; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_rs2_value <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_rs2_value <= issue_io_out_bits_0_rs2_value; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_imm <= issue_io_out_bits_0_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_rs1 <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_rs1 <= issue_io_out_bits_0_rs1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_dest <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_dest <= issue_io_out_bits_0_dest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_fu_type <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_fu_type <= issue_io_out_bits_0_fu_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_bru_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_bru_op <= issue_io_out_bits_0_bru_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_alu_op <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_alu_op <= issue_io_out_bits_0_alu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_lsu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_lsu_op <= issue_io_out_bits_0_lsu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_csr_op <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_csr_op <= issue_io_out_bits_0_csr_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_mdu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_mdu_op <= issue_io_out_bits_0_mdu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_wen <= issue_io_out_bits_0_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_rv64 <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_rv64 <= issue_io_out_bits_0_rv64; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_bp_br_taken <= issue_io_out_bits_0_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_bp_br_target <= issue_io_out_bits_0_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_0_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_0_bp_br_type <= issue_io_out_bits_0_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_valid <= issue_io_out_bits_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_pc <= issue_io_out_bits_1_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_inst <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_inst <= issue_io_out_bits_1_inst; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_src1_value <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_src1_value <= issue_io_out_bits_1_src1_value; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_src2_value <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_src2_value <= issue_io_out_bits_1_src2_value; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_rs2_value <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_rs2_value <= issue_io_out_bits_1_rs2_value; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_imm <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_imm <= issue_io_out_bits_1_imm; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_rs1 <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_rs1 <= issue_io_out_bits_1_rs1; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_dest <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_dest <= issue_io_out_bits_1_dest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_fu_type <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_fu_type <= issue_io_out_bits_1_fu_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_bru_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_bru_op <= issue_io_out_bits_1_bru_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_alu_op <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_alu_op <= issue_io_out_bits_1_alu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_lsu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_lsu_op <= issue_io_out_bits_1_lsu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_csr_op <= 3'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_csr_op <= issue_io_out_bits_1_csr_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_mdu_op <= 4'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_mdu_op <= issue_io_out_bits_1_mdu_op; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_wen <= issue_io_out_bits_1_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_rv64 <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_rv64 <= issue_io_out_bits_1_rv64; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_bp_br_taken <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_bp_br_taken <= issue_io_out_bits_1_bp_br_taken; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_bp_br_target <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_bp_br_target <= issue_io_out_bits_1_bp_br_target; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      exu_io_in_bits_r_1_bp_br_type <= 2'h0; // @[Reg.scala 27:20]
    end else if (fire_3) begin // @[Reg.scala 28:19]
      exu_io_in_bits_r_1_bp_br_type <= issue_io_out_bits_1_bp_br_type; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Connect.scala 6:24]
      valid_4 <= 1'h0; // @[Connect.scala 6:24]
    end else begin
      valid_4 <= _GEN_113;
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_0_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_0_valid <= exu_io_out_bits_0_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_0_pc <= 32'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_0_pc <= exu_io_out_bits_0_pc; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_0_final_result <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_0_final_result <= exu_io_out_bits_0_final_result; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_0_dest <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_0_dest <= exu_io_out_bits_0_dest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_0_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_0_wen <= exu_io_out_bits_0_wen; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_1_valid <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_1_valid <= exu_io_out_bits_1_valid; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_1_final_result <= 64'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_1_final_result <= exu_io_out_bits_1_final_result; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_1_dest <= 5'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_1_dest <= exu_io_out_bits_1_dest; // @[Reg.scala 28:23]
    end
    if (reset) begin // @[Reg.scala 27:20]
      wbu_io_in_bits_r_1_wen <= 1'h0; // @[Reg.scala 27:20]
    end else if (fire_4) begin // @[Reg.scala 28:19]
      wbu_io_in_bits_r_1_wen <= exu_io_out_bits_1_wen; // @[Reg.scala 28:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  iqueue_io_in_bits_r_pc = _RAND_1[31:0];
  _RAND_2 = {4{`RANDOM}};
  iqueue_io_in_bits_r_inst = _RAND_2[127:0];
  _RAND_3 = {1{`RANDOM}};
  iqueue_io_in_bits_r_uncache = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  iqueue_io_in_bits_r_offset = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  iqueue_io_in_bits_r_bp_br_offset = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  iqueue_io_in_bits_r_bp_br_taken = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  iqueue_io_in_bits_r_bp_br_target = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  iqueue_io_in_bits_r_bp_br_type = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  valid_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  idu_io_in_bits_r_0_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  idu_io_in_bits_r_0_pc = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  idu_io_in_bits_r_0_inst = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  idu_io_in_bits_r_0_bp_br_taken = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  idu_io_in_bits_r_0_bp_br_target = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  idu_io_in_bits_r_0_bp_br_type = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  idu_io_in_bits_r_1_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  idu_io_in_bits_r_1_pc = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  idu_io_in_bits_r_1_inst = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  idu_io_in_bits_r_1_bp_br_taken = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  idu_io_in_bits_r_1_bp_br_target = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  idu_io_in_bits_r_1_bp_br_type = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  valid_2 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  issue_io_in_bits_r_0_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  issue_io_in_bits_r_0_pc = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  issue_io_in_bits_r_0_inst = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  issue_io_in_bits_r_0_src1 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  issue_io_in_bits_r_0_src2 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  issue_io_in_bits_r_0_rs1 = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  issue_io_in_bits_r_0_rs2 = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  issue_io_in_bits_r_0_dest = _RAND_30[4:0];
  _RAND_31 = {2{`RANDOM}};
  issue_io_in_bits_r_0_imm = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  issue_io_in_bits_r_0_fu_type = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  issue_io_in_bits_r_0_bru_op = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  issue_io_in_bits_r_0_alu_op = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  issue_io_in_bits_r_0_lsu_op = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  issue_io_in_bits_r_0_csr_op = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  issue_io_in_bits_r_0_mdu_op = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  issue_io_in_bits_r_0_wen = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  issue_io_in_bits_r_0_rv64 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  issue_io_in_bits_r_0_bp_br_taken = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  issue_io_in_bits_r_0_bp_br_target = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  issue_io_in_bits_r_0_bp_br_type = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  issue_io_in_bits_r_1_valid = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  issue_io_in_bits_r_1_pc = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  issue_io_in_bits_r_1_inst = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  issue_io_in_bits_r_1_src1 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  issue_io_in_bits_r_1_src2 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  issue_io_in_bits_r_1_rs1 = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  issue_io_in_bits_r_1_rs2 = _RAND_49[4:0];
  _RAND_50 = {1{`RANDOM}};
  issue_io_in_bits_r_1_dest = _RAND_50[4:0];
  _RAND_51 = {2{`RANDOM}};
  issue_io_in_bits_r_1_imm = _RAND_51[63:0];
  _RAND_52 = {1{`RANDOM}};
  issue_io_in_bits_r_1_fu_type = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  issue_io_in_bits_r_1_bru_op = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  issue_io_in_bits_r_1_alu_op = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  issue_io_in_bits_r_1_lsu_op = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  issue_io_in_bits_r_1_csr_op = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  issue_io_in_bits_r_1_mdu_op = _RAND_57[3:0];
  _RAND_58 = {1{`RANDOM}};
  issue_io_in_bits_r_1_wen = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  issue_io_in_bits_r_1_rv64 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  issue_io_in_bits_r_1_bp_br_taken = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  issue_io_in_bits_r_1_bp_br_target = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  issue_io_in_bits_r_1_bp_br_type = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  valid_3 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  exu_io_in_bits_r_0_valid = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  exu_io_in_bits_r_0_pc = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  exu_io_in_bits_r_0_inst = _RAND_66[31:0];
  _RAND_67 = {2{`RANDOM}};
  exu_io_in_bits_r_0_src1_value = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  exu_io_in_bits_r_0_src2_value = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  exu_io_in_bits_r_0_rs2_value = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  exu_io_in_bits_r_0_imm = _RAND_70[63:0];
  _RAND_71 = {1{`RANDOM}};
  exu_io_in_bits_r_0_rs1 = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  exu_io_in_bits_r_0_dest = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  exu_io_in_bits_r_0_fu_type = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  exu_io_in_bits_r_0_bru_op = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  exu_io_in_bits_r_0_alu_op = _RAND_75[4:0];
  _RAND_76 = {1{`RANDOM}};
  exu_io_in_bits_r_0_lsu_op = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  exu_io_in_bits_r_0_csr_op = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  exu_io_in_bits_r_0_mdu_op = _RAND_78[3:0];
  _RAND_79 = {1{`RANDOM}};
  exu_io_in_bits_r_0_wen = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  exu_io_in_bits_r_0_rv64 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  exu_io_in_bits_r_0_bp_br_taken = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  exu_io_in_bits_r_0_bp_br_target = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  exu_io_in_bits_r_0_bp_br_type = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  exu_io_in_bits_r_1_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  exu_io_in_bits_r_1_pc = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  exu_io_in_bits_r_1_inst = _RAND_86[31:0];
  _RAND_87 = {2{`RANDOM}};
  exu_io_in_bits_r_1_src1_value = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  exu_io_in_bits_r_1_src2_value = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  exu_io_in_bits_r_1_rs2_value = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  exu_io_in_bits_r_1_imm = _RAND_90[63:0];
  _RAND_91 = {1{`RANDOM}};
  exu_io_in_bits_r_1_rs1 = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  exu_io_in_bits_r_1_dest = _RAND_92[4:0];
  _RAND_93 = {1{`RANDOM}};
  exu_io_in_bits_r_1_fu_type = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  exu_io_in_bits_r_1_bru_op = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  exu_io_in_bits_r_1_alu_op = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  exu_io_in_bits_r_1_lsu_op = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  exu_io_in_bits_r_1_csr_op = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  exu_io_in_bits_r_1_mdu_op = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  exu_io_in_bits_r_1_wen = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  exu_io_in_bits_r_1_rv64 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  exu_io_in_bits_r_1_bp_br_taken = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  exu_io_in_bits_r_1_bp_br_target = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  exu_io_in_bits_r_1_bp_br_type = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  valid_4 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  wbu_io_in_bits_r_0_valid = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  wbu_io_in_bits_r_0_pc = _RAND_106[31:0];
  _RAND_107 = {2{`RANDOM}};
  wbu_io_in_bits_r_0_final_result = _RAND_107[63:0];
  _RAND_108 = {1{`RANDOM}};
  wbu_io_in_bits_r_0_dest = _RAND_108[4:0];
  _RAND_109 = {1{`RANDOM}};
  wbu_io_in_bits_r_0_wen = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  wbu_io_in_bits_r_1_valid = _RAND_110[0:0];
  _RAND_111 = {2{`RANDOM}};
  wbu_io_in_bits_r_1_final_result = _RAND_111[63:0];
  _RAND_112 = {1{`RANDOM}};
  wbu_io_in_bits_r_1_dest = _RAND_112[4:0];
  _RAND_113 = {1{`RANDOM}};
  wbu_io_in_bits_r_1_wen = _RAND_113[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SramBridge(
  input          io_sram_cache_0_en,
  input          io_sram_cache_0_wen,
  input  [5:0]   io_sram_cache_0_addr,
  input  [127:0] io_sram_cache_0_wdata,
  output [127:0] io_sram_cache_0_rdata,
  input          io_sram_cache_1_en,
  input          io_sram_cache_1_wen,
  input  [5:0]   io_sram_cache_1_addr,
  input  [127:0] io_sram_cache_1_wdata,
  output [127:0] io_sram_cache_1_rdata,
  input          io_sram_cache_2_en,
  input          io_sram_cache_2_wen,
  input  [5:0]   io_sram_cache_2_addr,
  input  [127:0] io_sram_cache_2_wdata,
  output [127:0] io_sram_cache_2_rdata,
  input          io_sram_cache_3_en,
  input          io_sram_cache_3_wen,
  input  [5:0]   io_sram_cache_3_addr,
  input  [127:0] io_sram_cache_3_wdata,
  output [127:0] io_sram_cache_3_rdata,
  input          io_sram_cache_4_en,
  input          io_sram_cache_4_wen,
  input  [5:0]   io_sram_cache_4_addr,
  input  [127:0] io_sram_cache_4_wdata,
  output [127:0] io_sram_cache_4_rdata,
  input          io_sram_cache_5_en,
  input          io_sram_cache_5_wen,
  input  [5:0]   io_sram_cache_5_addr,
  input  [127:0] io_sram_cache_5_wdata,
  output [127:0] io_sram_cache_5_rdata,
  input          io_sram_cache_6_en,
  input          io_sram_cache_6_wen,
  input  [5:0]   io_sram_cache_6_addr,
  input  [127:0] io_sram_cache_6_wdata,
  output [127:0] io_sram_cache_6_rdata,
  input          io_sram_cache_7_en,
  input          io_sram_cache_7_wen,
  input  [5:0]   io_sram_cache_7_addr,
  input  [127:0] io_sram_cache_7_wdata,
  output [127:0] io_sram_cache_7_rdata,
  output [5:0]   io_sram_share_0_addr,
  output         io_sram_share_0_cen,
  output         io_sram_share_0_wen,
  output [127:0] io_sram_share_0_wdata,
  input  [127:0] io_sram_share_0_rdata,
  output [5:0]   io_sram_share_1_addr,
  output         io_sram_share_1_cen,
  output         io_sram_share_1_wen,
  output [127:0] io_sram_share_1_wdata,
  input  [127:0] io_sram_share_1_rdata,
  output [5:0]   io_sram_share_2_addr,
  output         io_sram_share_2_cen,
  output         io_sram_share_2_wen,
  output [127:0] io_sram_share_2_wdata,
  input  [127:0] io_sram_share_2_rdata,
  output [5:0]   io_sram_share_3_addr,
  output         io_sram_share_3_cen,
  output         io_sram_share_3_wen,
  output [127:0] io_sram_share_3_wdata,
  input  [127:0] io_sram_share_3_rdata,
  output [5:0]   io_sram_share_4_addr,
  output         io_sram_share_4_cen,
  output         io_sram_share_4_wen,
  output [127:0] io_sram_share_4_wdata,
  input  [127:0] io_sram_share_4_rdata,
  output [5:0]   io_sram_share_5_addr,
  output         io_sram_share_5_cen,
  output         io_sram_share_5_wen,
  output [127:0] io_sram_share_5_wdata,
  input  [127:0] io_sram_share_5_rdata,
  output [5:0]   io_sram_share_6_addr,
  output         io_sram_share_6_cen,
  output         io_sram_share_6_wen,
  output [127:0] io_sram_share_6_wdata,
  input  [127:0] io_sram_share_6_rdata,
  output [5:0]   io_sram_share_7_addr,
  output         io_sram_share_7_cen,
  output         io_sram_share_7_wen,
  output [127:0] io_sram_share_7_wdata,
  input  [127:0] io_sram_share_7_rdata
);
  assign io_sram_cache_0_rdata = io_sram_share_0_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_1_rdata = io_sram_share_1_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_2_rdata = io_sram_share_2_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_3_rdata = io_sram_share_3_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_4_rdata = io_sram_share_4_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_5_rdata = io_sram_share_5_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_6_rdata = io_sram_share_6_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_cache_7_rdata = io_sram_share_7_rdata; // @[SramBridge.scala 21:25]
  assign io_sram_share_0_addr = io_sram_cache_0_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_0_cen = ~io_sram_cache_0_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_0_wen = ~io_sram_cache_0_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_0_wdata = io_sram_cache_0_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_1_addr = io_sram_cache_1_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_1_cen = ~io_sram_cache_1_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_1_wen = ~io_sram_cache_1_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_1_wdata = io_sram_cache_1_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_2_addr = io_sram_cache_2_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_2_cen = ~io_sram_cache_2_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_2_wen = ~io_sram_cache_2_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_2_wdata = io_sram_cache_2_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_3_addr = io_sram_cache_3_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_3_cen = ~io_sram_cache_3_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_3_wen = ~io_sram_cache_3_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_3_wdata = io_sram_cache_3_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_4_addr = io_sram_cache_4_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_4_cen = ~io_sram_cache_4_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_4_wen = ~io_sram_cache_4_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_4_wdata = io_sram_cache_4_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_5_addr = io_sram_cache_5_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_5_cen = ~io_sram_cache_5_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_5_wen = ~io_sram_cache_5_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_5_wdata = io_sram_cache_5_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_6_addr = io_sram_cache_6_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_6_cen = ~io_sram_cache_6_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_6_wen = ~io_sram_cache_6_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_6_wdata = io_sram_cache_6_wdata; // @[SramBridge.scala 19:25]
  assign io_sram_share_7_addr = io_sram_cache_7_addr; // @[SramBridge.scala 15:24]
  assign io_sram_share_7_cen = ~io_sram_cache_7_en; // @[SramBridge.scala 16:26]
  assign io_sram_share_7_wen = ~io_sram_cache_7_wen; // @[SramBridge.scala 17:26]
  assign io_sram_share_7_wdata = io_sram_cache_7_wdata; // @[SramBridge.scala 19:25]
endmodule
module SocBridge(
  input          clock,
  input          reset,
  input          io_icache_rd_req,
  input  [2:0]   io_icache_rd_size,
  input  [31:0]  io_icache_rd_addr,
  output         io_icache_rd_rdy,
  output         io_icache_ret_valid,
  output [127:0] io_icache_ret_data,
  input          io_dcache_rd_req,
  input  [2:0]   io_dcache_rd_size,
  input  [31:0]  io_dcache_rd_addr,
  output         io_dcache_rd_rdy,
  output         io_dcache_ret_valid,
  output [127:0] io_dcache_ret_data,
  input          io_dcache_wr_req,
  input  [2:0]   io_dcache_wr_size,
  input  [31:0]  io_dcache_wr_addr,
  input  [7:0]   io_dcache_wr_wstrb,
  input  [127:0] io_dcache_wr_data,
  output         io_dcache_wr_rdy,
  output         io_dcache_wr_ok,
  input          io_out_awready,
  output         io_out_awvalid,
  output [31:0]  io_out_awaddr,
  output [7:0]   io_out_awlen,
  output [2:0]   io_out_awsize,
  input          io_out_wready,
  output         io_out_wvalid,
  output [63:0]  io_out_wdata,
  output [7:0]   io_out_wstrb,
  output         io_out_wlast,
  output         io_out_bready,
  input          io_out_bvalid,
  input          io_out_arready,
  output         io_out_arvalid,
  output [31:0]  io_out_araddr,
  output [3:0]   io_out_arid,
  output [7:0]   io_out_arlen,
  output [2:0]   io_out_arsize,
  output         io_out_rready,
  input          io_out_rvalid,
  input  [63:0]  io_out_rdata,
  input          io_out_rlast,
  input  [3:0]   io_out_rid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  ar_state; // @[SocBridge.scala 19:25]
  reg [1:0] w_state; // @[SocBridge.scala 20:24]
  reg  b_state; // @[SocBridge.scala 21:24]
  reg [3:0] arid; // @[SocBridge.scala 23:21]
  reg [31:0] araddr; // @[SocBridge.scala 24:23]
  reg [7:0] arlen; // @[SocBridge.scala 25:22]
  reg [2:0] arsize; // @[SocBridge.scala 26:23]
  reg [31:0] awaddr; // @[SocBridge.scala 28:23]
  reg [7:0] awlen; // @[SocBridge.scala 29:22]
  reg [2:0] awsize; // @[SocBridge.scala 30:23]
  reg [7:0] wstrb; // @[SocBridge.scala 31:22]
  reg [127:0] inst_rdata; // @[SocBridge.scala 33:27]
  reg [127:0] data_rdata; // @[SocBridge.scala 34:27]
  reg [127:0] data_wdata; // @[SocBridge.scala 35:27]
  reg  inst_rvalid; // @[SocBridge.scala 36:28]
  reg  data_rvalid; // @[SocBridge.scala 37:28]
  reg  wlast; // @[SocBridge.scala 38:22]
  wire [63:0] inst_rdata_lo = inst_rdata[63:0]; // @[SocBridge.scala 46:48]
  wire [127:0] _inst_rdata_T = {io_out_rdata,inst_rdata_lo}; // @[Cat.scala 30:58]
  wire [63:0] inst_rdata_hi = inst_rdata[127:64]; // @[SocBridge.scala 49:37]
  wire [127:0] _inst_rdata_T_1 = {inst_rdata_hi,io_out_rdata}; // @[Cat.scala 30:58]
  wire [63:0] data_rdata_lo = data_rdata[63:0]; // @[SocBridge.scala 53:48]
  wire [127:0] _data_rdata_T = {io_out_rdata,data_rdata_lo}; // @[Cat.scala 30:58]
  wire [63:0] data_rdata_hi = data_rdata[127:64]; // @[SocBridge.scala 56:37]
  wire [127:0] _data_rdata_T_1 = {data_rdata_hi,io_out_rdata}; // @[Cat.scala 30:58]
  wire  _GEN_4 = io_out_rid == 4'h0 & io_out_rlast; // @[SocBridge.scala 44:27 SocBridge.scala 40:15]
  wire  _GEN_6 = io_out_rid == 4'h0 ? 1'h0 : io_out_rlast; // @[SocBridge.scala 44:27 SocBridge.scala 41:15]
  wire  _GEN_8 = io_out_rvalid & io_out_rready & _GEN_4; // @[SocBridge.scala 43:34 SocBridge.scala 40:15]
  wire  _GEN_10 = io_out_rvalid & io_out_rready & _GEN_6; // @[SocBridge.scala 43:34 SocBridge.scala 41:15]
  wire  _T_2 = ~ar_state; // @[Conditional.scala 37:30]
  wire  _arlen_T_1 = io_dcache_rd_size == 3'h2 ? 1'h0 : 1'h1; // @[SocBridge.scala 67:21]
  wire  _arlen_T_3 = io_icache_rd_size == 3'h2 ? 1'h0 : 1'h1; // @[SocBridge.scala 73:21]
  wire  _GEN_11 = io_icache_rd_req & io_icache_rd_rdy | ar_state; // @[SocBridge.scala 69:50 SocBridge.scala 70:18 SocBridge.scala 19:25]
  wire  _GEN_16 = io_dcache_rd_req & io_dcache_rd_rdy | _GEN_11; // @[SocBridge.scala 63:44 SocBridge.scala 64:18]
  wire  _T_7 = 2'h0 == w_state; // @[Conditional.scala 37:30]
  wire  _awlen_T = io_dcache_wr_size == 3'h2; // @[SocBridge.scala 89:37]
  wire  _awlen_T_1 = io_dcache_wr_size == 3'h2 ? 1'h0 : 1'h1; // @[SocBridge.scala 89:21]
  wire  _T_9 = 2'h1 == w_state; // @[Conditional.scala 37:30]
  wire  _GEN_34 = awlen == 8'h0 | wlast; // @[SocBridge.scala 98:30 SocBridge.scala 99:17 SocBridge.scala 38:22]
  wire  _T_12 = 2'h2 == w_state; // @[Conditional.scala 37:30]
  wire  _T_13 = io_out_wvalid & io_out_wready; // @[SocBridge.scala 104:23]
  wire [1:0] _GEN_37 = _T_13 & wlast ? 2'h0 : w_state; // @[SocBridge.scala 107:53 SocBridge.scala 108:17 SocBridge.scala 20:24]
  wire  _GEN_38 = _T_13 & wlast ? 1'h0 : wlast; // @[SocBridge.scala 107:53 SocBridge.scala 109:15 SocBridge.scala 38:22]
  wire [1:0] _GEN_39 = io_out_wvalid & io_out_wready & ~wlast ? 2'h2 : _GEN_37; // @[SocBridge.scala 104:48 SocBridge.scala 105:17]
  wire  _GEN_40 = io_out_wvalid & io_out_wready & ~wlast | _GEN_38; // @[SocBridge.scala 104:48 SocBridge.scala 106:15]
  wire  _T_18 = ~b_state; // @[Conditional.scala 37:30]
  wire  _GEN_52 = io_out_bvalid & io_out_bready | b_state; // @[SocBridge.scala 116:38 SocBridge.scala 117:17 SocBridge.scala 21:24]
  assign io_icache_rd_rdy = _T_2 & ~io_dcache_rd_req; // @[SocBridge.scala 148:43]
  assign io_icache_ret_valid = inst_rvalid; // @[SocBridge.scala 149:20]
  assign io_icache_ret_data = inst_rdata; // @[SocBridge.scala 150:19]
  assign io_dcache_rd_rdy = ~ar_state; // @[SocBridge.scala 154:30]
  assign io_dcache_ret_valid = data_rvalid; // @[SocBridge.scala 155:20]
  assign io_dcache_ret_data = data_rdata; // @[SocBridge.scala 156:19]
  assign io_dcache_wr_rdy = w_state == 2'h0; // @[SocBridge.scala 157:29]
  assign io_dcache_wr_ok = b_state; // @[SocBridge.scala 158:28]
  assign io_out_awvalid = w_state == 2'h1; // @[SocBridge.scala 130:27]
  assign io_out_awaddr = awaddr; // @[SocBridge.scala 125:14]
  assign io_out_awlen = awlen; // @[SocBridge.scala 127:13]
  assign io_out_awsize = awsize; // @[SocBridge.scala 128:14]
  assign io_out_wvalid = w_state == 2'h2; // @[SocBridge.scala 135:26]
  assign io_out_wdata = wlast ? data_wdata[127:64] : data_wdata[63:0]; // @[SocBridge.scala 132:19]
  assign io_out_wstrb = wstrb; // @[SocBridge.scala 133:13]
  assign io_out_wlast = wlast; // @[SocBridge.scala 134:13]
  assign io_out_bready = ~b_state; // @[SocBridge.scala 146:26]
  assign io_out_arvalid = ar_state; // @[SocBridge.scala 142:28]
  assign io_out_araddr = araddr; // @[SocBridge.scala 137:14]
  assign io_out_arid = arid; // @[SocBridge.scala 138:12]
  assign io_out_arlen = arlen; // @[SocBridge.scala 139:13]
  assign io_out_arsize = arsize; // @[SocBridge.scala 140:14]
  assign io_out_rready = 1'h1; // @[SocBridge.scala 144:14]
  always @(posedge clock) begin
    if (reset) begin // @[SocBridge.scala 19:25]
      ar_state <= 1'h0; // @[SocBridge.scala 19:25]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      ar_state <= _GEN_16;
    end else if (ar_state) begin // @[Conditional.scala 39:67]
      if (io_out_arvalid & io_out_arready) begin // @[SocBridge.scala 78:40]
        ar_state <= 1'h0; // @[SocBridge.scala 79:18]
      end
    end
    if (reset) begin // @[SocBridge.scala 20:24]
      w_state <= 2'h0; // @[SocBridge.scala 20:24]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (io_dcache_wr_req & io_dcache_wr_rdy) begin // @[SocBridge.scala 86:44]
        w_state <= 2'h1; // @[SocBridge.scala 87:17]
      end
    end else if (_T_9) begin // @[Conditional.scala 39:67]
      if (io_out_awvalid & io_out_awready) begin // @[SocBridge.scala 96:40]
        w_state <= 2'h2; // @[SocBridge.scala 97:17]
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      w_state <= _GEN_39;
    end
    if (reset) begin // @[SocBridge.scala 21:24]
      b_state <= 1'h0; // @[SocBridge.scala 21:24]
    end else if (_T_18) begin // @[Conditional.scala 40:58]
      b_state <= _GEN_52;
    end else if (b_state) begin // @[Conditional.scala 39:67]
      b_state <= 1'h0; // @[SocBridge.scala 121:15]
    end
    if (reset) begin // @[SocBridge.scala 23:21]
      arid <= 4'h0; // @[SocBridge.scala 23:21]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_dcache_rd_req & io_dcache_rd_rdy) begin // @[SocBridge.scala 63:44]
        arid <= 4'h1; // @[SocBridge.scala 65:14]
      end else if (io_icache_rd_req & io_icache_rd_rdy) begin // @[SocBridge.scala 69:50]
        arid <= 4'h0; // @[SocBridge.scala 71:14]
      end
    end
    if (reset) begin // @[SocBridge.scala 24:23]
      araddr <= 32'h0; // @[SocBridge.scala 24:23]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_dcache_rd_req & io_dcache_rd_rdy) begin // @[SocBridge.scala 63:44]
        araddr <= io_dcache_rd_addr; // @[SocBridge.scala 66:16]
      end else if (io_icache_rd_req & io_icache_rd_rdy) begin // @[SocBridge.scala 69:50]
        araddr <= io_icache_rd_addr; // @[SocBridge.scala 72:16]
      end
    end
    if (reset) begin // @[SocBridge.scala 25:22]
      arlen <= 8'h0; // @[SocBridge.scala 25:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_dcache_rd_req & io_dcache_rd_rdy) begin // @[SocBridge.scala 63:44]
        arlen <= {{7'd0}, _arlen_T_1}; // @[SocBridge.scala 67:15]
      end else if (io_icache_rd_req & io_icache_rd_rdy) begin // @[SocBridge.scala 69:50]
        arlen <= {{7'd0}, _arlen_T_3}; // @[SocBridge.scala 73:15]
      end
    end
    if (reset) begin // @[SocBridge.scala 26:23]
      arsize <= 3'h0; // @[SocBridge.scala 26:23]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io_dcache_rd_req & io_dcache_rd_rdy) begin // @[SocBridge.scala 63:44]
        arsize <= io_dcache_rd_size; // @[SocBridge.scala 68:16]
      end else if (io_icache_rd_req & io_icache_rd_rdy) begin // @[SocBridge.scala 69:50]
        arsize <= io_icache_rd_size; // @[SocBridge.scala 74:16]
      end
    end
    if (reset) begin // @[SocBridge.scala 28:23]
      awaddr <= 32'h0; // @[SocBridge.scala 28:23]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (io_dcache_wr_req & io_dcache_wr_rdy) begin // @[SocBridge.scala 86:44]
        awaddr <= io_dcache_wr_addr; // @[SocBridge.scala 88:16]
      end
    end
    if (reset) begin // @[SocBridge.scala 29:22]
      awlen <= 8'h0; // @[SocBridge.scala 29:22]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (io_dcache_wr_req & io_dcache_wr_rdy) begin // @[SocBridge.scala 86:44]
        awlen <= {{7'd0}, _awlen_T_1}; // @[SocBridge.scala 89:15]
      end
    end
    if (reset) begin // @[SocBridge.scala 30:23]
      awsize <= 3'h0; // @[SocBridge.scala 30:23]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (io_dcache_wr_req & io_dcache_wr_rdy) begin // @[SocBridge.scala 86:44]
        awsize <= io_dcache_wr_size; // @[SocBridge.scala 90:16]
      end
    end
    if (reset) begin // @[SocBridge.scala 31:22]
      wstrb <= 8'h0; // @[SocBridge.scala 31:22]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (io_dcache_wr_req & io_dcache_wr_rdy) begin // @[SocBridge.scala 86:44]
        if (_awlen_T) begin // @[SocBridge.scala 91:21]
          wstrb <= io_dcache_wr_wstrb;
        end else begin
          wstrb <= 8'hff;
        end
      end
    end
    if (reset) begin // @[SocBridge.scala 33:27]
      inst_rdata <= 128'h0; // @[SocBridge.scala 33:27]
    end else if (io_out_rvalid & io_out_rready) begin // @[SocBridge.scala 43:34]
      if (io_out_rid == 4'h0) begin // @[SocBridge.scala 44:27]
        if (io_out_rlast) begin // @[SocBridge.scala 45:23]
          inst_rdata <= _inst_rdata_T; // @[SocBridge.scala 46:20]
        end else begin
          inst_rdata <= _inst_rdata_T_1; // @[SocBridge.scala 49:20]
        end
      end
    end
    if (reset) begin // @[SocBridge.scala 34:27]
      data_rdata <= 128'h0; // @[SocBridge.scala 34:27]
    end else if (io_out_rvalid & io_out_rready) begin // @[SocBridge.scala 43:34]
      if (!(io_out_rid == 4'h0)) begin // @[SocBridge.scala 44:27]
        if (io_out_rlast) begin // @[SocBridge.scala 52:23]
          data_rdata <= _data_rdata_T; // @[SocBridge.scala 53:20]
        end else begin
          data_rdata <= _data_rdata_T_1; // @[SocBridge.scala 56:20]
        end
      end
    end
    if (reset) begin // @[SocBridge.scala 35:27]
      data_wdata <= 128'h0; // @[SocBridge.scala 35:27]
    end else if (_T_7) begin // @[Conditional.scala 40:58]
      if (io_dcache_wr_req & io_dcache_wr_rdy) begin // @[SocBridge.scala 86:44]
        data_wdata <= io_dcache_wr_data; // @[SocBridge.scala 92:20]
      end
    end
    if (reset) begin // @[SocBridge.scala 36:28]
      inst_rvalid <= 1'h0; // @[SocBridge.scala 36:28]
    end else begin
      inst_rvalid <= _GEN_8;
    end
    if (reset) begin // @[SocBridge.scala 37:28]
      data_rvalid <= 1'h0; // @[SocBridge.scala 37:28]
    end else begin
      data_rvalid <= _GEN_10;
    end
    if (reset) begin // @[SocBridge.scala 38:22]
      wlast <= 1'h0; // @[SocBridge.scala 38:22]
    end else if (!(_T_7)) begin // @[Conditional.scala 40:58]
      if (_T_9) begin // @[Conditional.scala 39:67]
        if (io_out_awvalid & io_out_awready) begin // @[SocBridge.scala 96:40]
          wlast <= _GEN_34;
        end
      end else if (_T_12) begin // @[Conditional.scala 39:67]
        wlast <= _GEN_40;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  w_state = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  b_state = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  arid = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  araddr = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  arlen = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  arsize = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  awaddr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  awlen = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  awsize = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  wstrb = _RAND_10[7:0];
  _RAND_11 = {4{`RANDOM}};
  inst_rdata = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  data_rdata = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  data_wdata = _RAND_13[127:0];
  _RAND_14 = {1{`RANDOM}};
  inst_rvalid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  data_rvalid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  wlast = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SocTop(
  input          clock,
  input          reset,
  input          io_master_awready,
  output         io_master_awvalid,
  output [31:0]  io_master_awaddr,
  output [7:0]   io_master_awlen,
  output [2:0]   io_master_awsize,
  input          io_master_wready,
  output         io_master_wvalid,
  output [63:0]  io_master_wdata,
  output [7:0]   io_master_wstrb,
  output         io_master_wlast,
  output         io_master_bready,
  input          io_master_bvalid,
  input          io_master_arready,
  output         io_master_arvalid,
  output [31:0]  io_master_araddr,
  output [3:0]   io_master_arid,
  output [7:0]   io_master_arlen,
  output [2:0]   io_master_arsize,
  input          io_master_rvalid,
  input  [63:0]  io_master_rdata,
  input          io_master_rlast,
  input  [3:0]   io_master_rid,
  output [5:0]   io_sram0_addr,
  output         io_sram0_cen,
  output         io_sram0_wen,
  output [127:0] io_sram0_wdata,
  input  [127:0] io_sram0_rdata,
  output [5:0]   io_sram1_addr,
  output         io_sram1_cen,
  output         io_sram1_wen,
  output [127:0] io_sram1_wdata,
  input  [127:0] io_sram1_rdata,
  output [5:0]   io_sram2_addr,
  output         io_sram2_cen,
  output         io_sram2_wen,
  output [127:0] io_sram2_wdata,
  input  [127:0] io_sram2_rdata,
  output [5:0]   io_sram3_addr,
  output         io_sram3_cen,
  output         io_sram3_wen,
  output [127:0] io_sram3_wdata,
  input  [127:0] io_sram3_rdata,
  output [5:0]   io_sram4_addr,
  output         io_sram4_cen,
  output         io_sram4_wen,
  output [127:0] io_sram4_wdata,
  input  [127:0] io_sram4_rdata,
  output [5:0]   io_sram5_addr,
  output         io_sram5_cen,
  output         io_sram5_wen,
  output [127:0] io_sram5_wdata,
  input  [127:0] io_sram5_rdata,
  output [5:0]   io_sram6_addr,
  output         io_sram6_cen,
  output         io_sram6_wen,
  output [127:0] io_sram6_wdata,
  input  [127:0] io_sram6_rdata,
  output [5:0]   io_sram7_addr,
  output         io_sram7_cen,
  output         io_sram7_wen,
  output [127:0] io_sram7_wdata,
  input  [127:0] io_sram7_rdata,
  output [31:0]  io_commit_0_pc
);
  wire  core_clock; // @[SocTop.scala 19:20]
  wire  core_reset; // @[SocTop.scala 19:20]
  wire  core_io_icache_bridge_rd_req; // @[SocTop.scala 19:20]
  wire [2:0] core_io_icache_bridge_rd_size; // @[SocTop.scala 19:20]
  wire [31:0] core_io_icache_bridge_rd_addr; // @[SocTop.scala 19:20]
  wire  core_io_icache_bridge_rd_rdy; // @[SocTop.scala 19:20]
  wire  core_io_icache_bridge_ret_valid; // @[SocTop.scala 19:20]
  wire [127:0] core_io_icache_bridge_ret_data; // @[SocTop.scala 19:20]
  wire  core_io_dcache_bridge_rd_req; // @[SocTop.scala 19:20]
  wire [2:0] core_io_dcache_bridge_rd_size; // @[SocTop.scala 19:20]
  wire [31:0] core_io_dcache_bridge_rd_addr; // @[SocTop.scala 19:20]
  wire  core_io_dcache_bridge_rd_rdy; // @[SocTop.scala 19:20]
  wire  core_io_dcache_bridge_ret_valid; // @[SocTop.scala 19:20]
  wire [127:0] core_io_dcache_bridge_ret_data; // @[SocTop.scala 19:20]
  wire  core_io_dcache_bridge_wr_req; // @[SocTop.scala 19:20]
  wire [2:0] core_io_dcache_bridge_wr_size; // @[SocTop.scala 19:20]
  wire [31:0] core_io_dcache_bridge_wr_addr; // @[SocTop.scala 19:20]
  wire [7:0] core_io_dcache_bridge_wr_wstrb; // @[SocTop.scala 19:20]
  wire [127:0] core_io_dcache_bridge_wr_data; // @[SocTop.scala 19:20]
  wire  core_io_dcache_bridge_wr_rdy; // @[SocTop.scala 19:20]
  wire  core_io_dcache_bridge_wr_ok; // @[SocTop.scala 19:20]
  wire  core_io_sram_0_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_0_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_0_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_0_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_0_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_1_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_1_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_1_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_1_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_1_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_2_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_2_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_2_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_2_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_2_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_3_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_3_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_3_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_3_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_3_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_4_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_4_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_4_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_4_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_4_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_5_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_5_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_5_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_5_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_5_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_6_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_6_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_6_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_6_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_6_rdata; // @[SocTop.scala 19:20]
  wire  core_io_sram_7_en; // @[SocTop.scala 19:20]
  wire  core_io_sram_7_wen; // @[SocTop.scala 19:20]
  wire [5:0] core_io_sram_7_addr; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_7_wdata; // @[SocTop.scala 19:20]
  wire [127:0] core_io_sram_7_rdata; // @[SocTop.scala 19:20]
  wire [31:0] core_io_commit_0_pc; // @[SocTop.scala 19:20]
  wire  sram_bridge_io_sram_cache_0_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_0_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_0_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_0_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_0_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_1_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_1_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_1_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_1_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_1_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_2_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_2_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_2_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_2_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_2_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_3_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_3_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_3_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_3_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_3_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_4_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_4_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_4_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_4_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_4_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_5_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_5_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_5_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_5_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_5_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_6_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_6_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_6_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_6_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_6_rdata; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_7_en; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_cache_7_wen; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_cache_7_addr; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_7_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_cache_7_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_0_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_0_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_0_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_0_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_0_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_1_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_1_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_1_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_1_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_1_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_2_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_2_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_2_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_2_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_2_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_3_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_3_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_3_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_3_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_3_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_4_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_4_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_4_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_4_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_4_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_5_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_5_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_5_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_5_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_5_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_6_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_6_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_6_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_6_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_6_rdata; // @[SocTop.scala 20:27]
  wire [5:0] sram_bridge_io_sram_share_7_addr; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_7_cen; // @[SocTop.scala 20:27]
  wire  sram_bridge_io_sram_share_7_wen; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_7_wdata; // @[SocTop.scala 20:27]
  wire [127:0] sram_bridge_io_sram_share_7_rdata; // @[SocTop.scala 20:27]
  wire  transfer_bridge_clock; // @[SocTop.scala 31:31]
  wire  transfer_bridge_reset; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_icache_rd_req; // @[SocTop.scala 31:31]
  wire [2:0] transfer_bridge_io_icache_rd_size; // @[SocTop.scala 31:31]
  wire [31:0] transfer_bridge_io_icache_rd_addr; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_icache_rd_rdy; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_icache_ret_valid; // @[SocTop.scala 31:31]
  wire [127:0] transfer_bridge_io_icache_ret_data; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_dcache_rd_req; // @[SocTop.scala 31:31]
  wire [2:0] transfer_bridge_io_dcache_rd_size; // @[SocTop.scala 31:31]
  wire [31:0] transfer_bridge_io_dcache_rd_addr; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_dcache_rd_rdy; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_dcache_ret_valid; // @[SocTop.scala 31:31]
  wire [127:0] transfer_bridge_io_dcache_ret_data; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_dcache_wr_req; // @[SocTop.scala 31:31]
  wire [2:0] transfer_bridge_io_dcache_wr_size; // @[SocTop.scala 31:31]
  wire [31:0] transfer_bridge_io_dcache_wr_addr; // @[SocTop.scala 31:31]
  wire [7:0] transfer_bridge_io_dcache_wr_wstrb; // @[SocTop.scala 31:31]
  wire [127:0] transfer_bridge_io_dcache_wr_data; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_dcache_wr_rdy; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_dcache_wr_ok; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_awready; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_awvalid; // @[SocTop.scala 31:31]
  wire [31:0] transfer_bridge_io_out_awaddr; // @[SocTop.scala 31:31]
  wire [7:0] transfer_bridge_io_out_awlen; // @[SocTop.scala 31:31]
  wire [2:0] transfer_bridge_io_out_awsize; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_wready; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_wvalid; // @[SocTop.scala 31:31]
  wire [63:0] transfer_bridge_io_out_wdata; // @[SocTop.scala 31:31]
  wire [7:0] transfer_bridge_io_out_wstrb; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_wlast; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_bready; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_bvalid; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_arready; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_arvalid; // @[SocTop.scala 31:31]
  wire [31:0] transfer_bridge_io_out_araddr; // @[SocTop.scala 31:31]
  wire [3:0] transfer_bridge_io_out_arid; // @[SocTop.scala 31:31]
  wire [7:0] transfer_bridge_io_out_arlen; // @[SocTop.scala 31:31]
  wire [2:0] transfer_bridge_io_out_arsize; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_rready; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_rvalid; // @[SocTop.scala 31:31]
  wire [63:0] transfer_bridge_io_out_rdata; // @[SocTop.scala 31:31]
  wire  transfer_bridge_io_out_rlast; // @[SocTop.scala 31:31]
  wire [3:0] transfer_bridge_io_out_rid; // @[SocTop.scala 31:31]
  Core_Soc core ( // @[SocTop.scala 19:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_icache_bridge_rd_req(core_io_icache_bridge_rd_req),
    .io_icache_bridge_rd_size(core_io_icache_bridge_rd_size),
    .io_icache_bridge_rd_addr(core_io_icache_bridge_rd_addr),
    .io_icache_bridge_rd_rdy(core_io_icache_bridge_rd_rdy),
    .io_icache_bridge_ret_valid(core_io_icache_bridge_ret_valid),
    .io_icache_bridge_ret_data(core_io_icache_bridge_ret_data),
    .io_dcache_bridge_rd_req(core_io_dcache_bridge_rd_req),
    .io_dcache_bridge_rd_size(core_io_dcache_bridge_rd_size),
    .io_dcache_bridge_rd_addr(core_io_dcache_bridge_rd_addr),
    .io_dcache_bridge_rd_rdy(core_io_dcache_bridge_rd_rdy),
    .io_dcache_bridge_ret_valid(core_io_dcache_bridge_ret_valid),
    .io_dcache_bridge_ret_data(core_io_dcache_bridge_ret_data),
    .io_dcache_bridge_wr_req(core_io_dcache_bridge_wr_req),
    .io_dcache_bridge_wr_size(core_io_dcache_bridge_wr_size),
    .io_dcache_bridge_wr_addr(core_io_dcache_bridge_wr_addr),
    .io_dcache_bridge_wr_wstrb(core_io_dcache_bridge_wr_wstrb),
    .io_dcache_bridge_wr_data(core_io_dcache_bridge_wr_data),
    .io_dcache_bridge_wr_rdy(core_io_dcache_bridge_wr_rdy),
    .io_dcache_bridge_wr_ok(core_io_dcache_bridge_wr_ok),
    .io_sram_0_en(core_io_sram_0_en),
    .io_sram_0_wen(core_io_sram_0_wen),
    .io_sram_0_addr(core_io_sram_0_addr),
    .io_sram_0_wdata(core_io_sram_0_wdata),
    .io_sram_0_rdata(core_io_sram_0_rdata),
    .io_sram_1_en(core_io_sram_1_en),
    .io_sram_1_wen(core_io_sram_1_wen),
    .io_sram_1_addr(core_io_sram_1_addr),
    .io_sram_1_wdata(core_io_sram_1_wdata),
    .io_sram_1_rdata(core_io_sram_1_rdata),
    .io_sram_2_en(core_io_sram_2_en),
    .io_sram_2_wen(core_io_sram_2_wen),
    .io_sram_2_addr(core_io_sram_2_addr),
    .io_sram_2_wdata(core_io_sram_2_wdata),
    .io_sram_2_rdata(core_io_sram_2_rdata),
    .io_sram_3_en(core_io_sram_3_en),
    .io_sram_3_wen(core_io_sram_3_wen),
    .io_sram_3_addr(core_io_sram_3_addr),
    .io_sram_3_wdata(core_io_sram_3_wdata),
    .io_sram_3_rdata(core_io_sram_3_rdata),
    .io_sram_4_en(core_io_sram_4_en),
    .io_sram_4_wen(core_io_sram_4_wen),
    .io_sram_4_addr(core_io_sram_4_addr),
    .io_sram_4_wdata(core_io_sram_4_wdata),
    .io_sram_4_rdata(core_io_sram_4_rdata),
    .io_sram_5_en(core_io_sram_5_en),
    .io_sram_5_wen(core_io_sram_5_wen),
    .io_sram_5_addr(core_io_sram_5_addr),
    .io_sram_5_wdata(core_io_sram_5_wdata),
    .io_sram_5_rdata(core_io_sram_5_rdata),
    .io_sram_6_en(core_io_sram_6_en),
    .io_sram_6_wen(core_io_sram_6_wen),
    .io_sram_6_addr(core_io_sram_6_addr),
    .io_sram_6_wdata(core_io_sram_6_wdata),
    .io_sram_6_rdata(core_io_sram_6_rdata),
    .io_sram_7_en(core_io_sram_7_en),
    .io_sram_7_wen(core_io_sram_7_wen),
    .io_sram_7_addr(core_io_sram_7_addr),
    .io_sram_7_wdata(core_io_sram_7_wdata),
    .io_sram_7_rdata(core_io_sram_7_rdata),
    .io_commit_0_pc(core_io_commit_0_pc)
  );
  SramBridge sram_bridge ( // @[SocTop.scala 20:27]
    .io_sram_cache_0_en(sram_bridge_io_sram_cache_0_en),
    .io_sram_cache_0_wen(sram_bridge_io_sram_cache_0_wen),
    .io_sram_cache_0_addr(sram_bridge_io_sram_cache_0_addr),
    .io_sram_cache_0_wdata(sram_bridge_io_sram_cache_0_wdata),
    .io_sram_cache_0_rdata(sram_bridge_io_sram_cache_0_rdata),
    .io_sram_cache_1_en(sram_bridge_io_sram_cache_1_en),
    .io_sram_cache_1_wen(sram_bridge_io_sram_cache_1_wen),
    .io_sram_cache_1_addr(sram_bridge_io_sram_cache_1_addr),
    .io_sram_cache_1_wdata(sram_bridge_io_sram_cache_1_wdata),
    .io_sram_cache_1_rdata(sram_bridge_io_sram_cache_1_rdata),
    .io_sram_cache_2_en(sram_bridge_io_sram_cache_2_en),
    .io_sram_cache_2_wen(sram_bridge_io_sram_cache_2_wen),
    .io_sram_cache_2_addr(sram_bridge_io_sram_cache_2_addr),
    .io_sram_cache_2_wdata(sram_bridge_io_sram_cache_2_wdata),
    .io_sram_cache_2_rdata(sram_bridge_io_sram_cache_2_rdata),
    .io_sram_cache_3_en(sram_bridge_io_sram_cache_3_en),
    .io_sram_cache_3_wen(sram_bridge_io_sram_cache_3_wen),
    .io_sram_cache_3_addr(sram_bridge_io_sram_cache_3_addr),
    .io_sram_cache_3_wdata(sram_bridge_io_sram_cache_3_wdata),
    .io_sram_cache_3_rdata(sram_bridge_io_sram_cache_3_rdata),
    .io_sram_cache_4_en(sram_bridge_io_sram_cache_4_en),
    .io_sram_cache_4_wen(sram_bridge_io_sram_cache_4_wen),
    .io_sram_cache_4_addr(sram_bridge_io_sram_cache_4_addr),
    .io_sram_cache_4_wdata(sram_bridge_io_sram_cache_4_wdata),
    .io_sram_cache_4_rdata(sram_bridge_io_sram_cache_4_rdata),
    .io_sram_cache_5_en(sram_bridge_io_sram_cache_5_en),
    .io_sram_cache_5_wen(sram_bridge_io_sram_cache_5_wen),
    .io_sram_cache_5_addr(sram_bridge_io_sram_cache_5_addr),
    .io_sram_cache_5_wdata(sram_bridge_io_sram_cache_5_wdata),
    .io_sram_cache_5_rdata(sram_bridge_io_sram_cache_5_rdata),
    .io_sram_cache_6_en(sram_bridge_io_sram_cache_6_en),
    .io_sram_cache_6_wen(sram_bridge_io_sram_cache_6_wen),
    .io_sram_cache_6_addr(sram_bridge_io_sram_cache_6_addr),
    .io_sram_cache_6_wdata(sram_bridge_io_sram_cache_6_wdata),
    .io_sram_cache_6_rdata(sram_bridge_io_sram_cache_6_rdata),
    .io_sram_cache_7_en(sram_bridge_io_sram_cache_7_en),
    .io_sram_cache_7_wen(sram_bridge_io_sram_cache_7_wen),
    .io_sram_cache_7_addr(sram_bridge_io_sram_cache_7_addr),
    .io_sram_cache_7_wdata(sram_bridge_io_sram_cache_7_wdata),
    .io_sram_cache_7_rdata(sram_bridge_io_sram_cache_7_rdata),
    .io_sram_share_0_addr(sram_bridge_io_sram_share_0_addr),
    .io_sram_share_0_cen(sram_bridge_io_sram_share_0_cen),
    .io_sram_share_0_wen(sram_bridge_io_sram_share_0_wen),
    .io_sram_share_0_wdata(sram_bridge_io_sram_share_0_wdata),
    .io_sram_share_0_rdata(sram_bridge_io_sram_share_0_rdata),
    .io_sram_share_1_addr(sram_bridge_io_sram_share_1_addr),
    .io_sram_share_1_cen(sram_bridge_io_sram_share_1_cen),
    .io_sram_share_1_wen(sram_bridge_io_sram_share_1_wen),
    .io_sram_share_1_wdata(sram_bridge_io_sram_share_1_wdata),
    .io_sram_share_1_rdata(sram_bridge_io_sram_share_1_rdata),
    .io_sram_share_2_addr(sram_bridge_io_sram_share_2_addr),
    .io_sram_share_2_cen(sram_bridge_io_sram_share_2_cen),
    .io_sram_share_2_wen(sram_bridge_io_sram_share_2_wen),
    .io_sram_share_2_wdata(sram_bridge_io_sram_share_2_wdata),
    .io_sram_share_2_rdata(sram_bridge_io_sram_share_2_rdata),
    .io_sram_share_3_addr(sram_bridge_io_sram_share_3_addr),
    .io_sram_share_3_cen(sram_bridge_io_sram_share_3_cen),
    .io_sram_share_3_wen(sram_bridge_io_sram_share_3_wen),
    .io_sram_share_3_wdata(sram_bridge_io_sram_share_3_wdata),
    .io_sram_share_3_rdata(sram_bridge_io_sram_share_3_rdata),
    .io_sram_share_4_addr(sram_bridge_io_sram_share_4_addr),
    .io_sram_share_4_cen(sram_bridge_io_sram_share_4_cen),
    .io_sram_share_4_wen(sram_bridge_io_sram_share_4_wen),
    .io_sram_share_4_wdata(sram_bridge_io_sram_share_4_wdata),
    .io_sram_share_4_rdata(sram_bridge_io_sram_share_4_rdata),
    .io_sram_share_5_addr(sram_bridge_io_sram_share_5_addr),
    .io_sram_share_5_cen(sram_bridge_io_sram_share_5_cen),
    .io_sram_share_5_wen(sram_bridge_io_sram_share_5_wen),
    .io_sram_share_5_wdata(sram_bridge_io_sram_share_5_wdata),
    .io_sram_share_5_rdata(sram_bridge_io_sram_share_5_rdata),
    .io_sram_share_6_addr(sram_bridge_io_sram_share_6_addr),
    .io_sram_share_6_cen(sram_bridge_io_sram_share_6_cen),
    .io_sram_share_6_wen(sram_bridge_io_sram_share_6_wen),
    .io_sram_share_6_wdata(sram_bridge_io_sram_share_6_wdata),
    .io_sram_share_6_rdata(sram_bridge_io_sram_share_6_rdata),
    .io_sram_share_7_addr(sram_bridge_io_sram_share_7_addr),
    .io_sram_share_7_cen(sram_bridge_io_sram_share_7_cen),
    .io_sram_share_7_wen(sram_bridge_io_sram_share_7_wen),
    .io_sram_share_7_wdata(sram_bridge_io_sram_share_7_wdata),
    .io_sram_share_7_rdata(sram_bridge_io_sram_share_7_rdata)
  );
  SocBridge transfer_bridge ( // @[SocTop.scala 31:31]
    .clock(transfer_bridge_clock),
    .reset(transfer_bridge_reset),
    .io_icache_rd_req(transfer_bridge_io_icache_rd_req),
    .io_icache_rd_size(transfer_bridge_io_icache_rd_size),
    .io_icache_rd_addr(transfer_bridge_io_icache_rd_addr),
    .io_icache_rd_rdy(transfer_bridge_io_icache_rd_rdy),
    .io_icache_ret_valid(transfer_bridge_io_icache_ret_valid),
    .io_icache_ret_data(transfer_bridge_io_icache_ret_data),
    .io_dcache_rd_req(transfer_bridge_io_dcache_rd_req),
    .io_dcache_rd_size(transfer_bridge_io_dcache_rd_size),
    .io_dcache_rd_addr(transfer_bridge_io_dcache_rd_addr),
    .io_dcache_rd_rdy(transfer_bridge_io_dcache_rd_rdy),
    .io_dcache_ret_valid(transfer_bridge_io_dcache_ret_valid),
    .io_dcache_ret_data(transfer_bridge_io_dcache_ret_data),
    .io_dcache_wr_req(transfer_bridge_io_dcache_wr_req),
    .io_dcache_wr_size(transfer_bridge_io_dcache_wr_size),
    .io_dcache_wr_addr(transfer_bridge_io_dcache_wr_addr),
    .io_dcache_wr_wstrb(transfer_bridge_io_dcache_wr_wstrb),
    .io_dcache_wr_data(transfer_bridge_io_dcache_wr_data),
    .io_dcache_wr_rdy(transfer_bridge_io_dcache_wr_rdy),
    .io_dcache_wr_ok(transfer_bridge_io_dcache_wr_ok),
    .io_out_awready(transfer_bridge_io_out_awready),
    .io_out_awvalid(transfer_bridge_io_out_awvalid),
    .io_out_awaddr(transfer_bridge_io_out_awaddr),
    .io_out_awlen(transfer_bridge_io_out_awlen),
    .io_out_awsize(transfer_bridge_io_out_awsize),
    .io_out_wready(transfer_bridge_io_out_wready),
    .io_out_wvalid(transfer_bridge_io_out_wvalid),
    .io_out_wdata(transfer_bridge_io_out_wdata),
    .io_out_wstrb(transfer_bridge_io_out_wstrb),
    .io_out_wlast(transfer_bridge_io_out_wlast),
    .io_out_bready(transfer_bridge_io_out_bready),
    .io_out_bvalid(transfer_bridge_io_out_bvalid),
    .io_out_arready(transfer_bridge_io_out_arready),
    .io_out_arvalid(transfer_bridge_io_out_arvalid),
    .io_out_araddr(transfer_bridge_io_out_araddr),
    .io_out_arid(transfer_bridge_io_out_arid),
    .io_out_arlen(transfer_bridge_io_out_arlen),
    .io_out_arsize(transfer_bridge_io_out_arsize),
    .io_out_rready(transfer_bridge_io_out_rready),
    .io_out_rvalid(transfer_bridge_io_out_rvalid),
    .io_out_rdata(transfer_bridge_io_out_rdata),
    .io_out_rlast(transfer_bridge_io_out_rlast),
    .io_out_rid(transfer_bridge_io_out_rid)
  );
  assign io_master_awvalid = transfer_bridge_io_out_awvalid; // @[SocTop.scala 34:26]
  assign io_master_awaddr = transfer_bridge_io_out_awaddr; // @[SocTop.scala 34:26]
  assign io_master_awlen = transfer_bridge_io_out_awlen; // @[SocTop.scala 34:26]
  assign io_master_awsize = transfer_bridge_io_out_awsize; // @[SocTop.scala 34:26]
  assign io_master_wvalid = transfer_bridge_io_out_wvalid; // @[SocTop.scala 34:26]
  assign io_master_wdata = transfer_bridge_io_out_wdata; // @[SocTop.scala 34:26]
  assign io_master_wstrb = transfer_bridge_io_out_wstrb; // @[SocTop.scala 34:26]
  assign io_master_wlast = transfer_bridge_io_out_wlast; // @[SocTop.scala 34:26]
  assign io_master_bready = transfer_bridge_io_out_bready; // @[SocTop.scala 34:26]
  assign io_master_arvalid = transfer_bridge_io_out_arvalid; // @[SocTop.scala 34:26]
  assign io_master_araddr = transfer_bridge_io_out_araddr; // @[SocTop.scala 34:26]
  assign io_master_arid = transfer_bridge_io_out_arid; // @[SocTop.scala 34:26]
  assign io_master_arlen = transfer_bridge_io_out_arlen; // @[SocTop.scala 34:26]
  assign io_master_arsize = transfer_bridge_io_out_arsize; // @[SocTop.scala 34:26]
  assign io_sram0_addr = sram_bridge_io_sram_share_0_addr; // @[SocTop.scala 22:32]
  assign io_sram0_cen = sram_bridge_io_sram_share_0_cen; // @[SocTop.scala 22:32]
  assign io_sram0_wen = sram_bridge_io_sram_share_0_wen; // @[SocTop.scala 22:32]
  assign io_sram0_wdata = sram_bridge_io_sram_share_0_wdata; // @[SocTop.scala 22:32]
  assign io_sram1_addr = sram_bridge_io_sram_share_1_addr; // @[SocTop.scala 23:32]
  assign io_sram1_cen = sram_bridge_io_sram_share_1_cen; // @[SocTop.scala 23:32]
  assign io_sram1_wen = sram_bridge_io_sram_share_1_wen; // @[SocTop.scala 23:32]
  assign io_sram1_wdata = sram_bridge_io_sram_share_1_wdata; // @[SocTop.scala 23:32]
  assign io_sram2_addr = sram_bridge_io_sram_share_2_addr; // @[SocTop.scala 24:32]
  assign io_sram2_cen = sram_bridge_io_sram_share_2_cen; // @[SocTop.scala 24:32]
  assign io_sram2_wen = sram_bridge_io_sram_share_2_wen; // @[SocTop.scala 24:32]
  assign io_sram2_wdata = sram_bridge_io_sram_share_2_wdata; // @[SocTop.scala 24:32]
  assign io_sram3_addr = sram_bridge_io_sram_share_3_addr; // @[SocTop.scala 25:32]
  assign io_sram3_cen = sram_bridge_io_sram_share_3_cen; // @[SocTop.scala 25:32]
  assign io_sram3_wen = sram_bridge_io_sram_share_3_wen; // @[SocTop.scala 25:32]
  assign io_sram3_wdata = sram_bridge_io_sram_share_3_wdata; // @[SocTop.scala 25:32]
  assign io_sram4_addr = sram_bridge_io_sram_share_4_addr; // @[SocTop.scala 26:32]
  assign io_sram4_cen = sram_bridge_io_sram_share_4_cen; // @[SocTop.scala 26:32]
  assign io_sram4_wen = sram_bridge_io_sram_share_4_wen; // @[SocTop.scala 26:32]
  assign io_sram4_wdata = sram_bridge_io_sram_share_4_wdata; // @[SocTop.scala 26:32]
  assign io_sram5_addr = sram_bridge_io_sram_share_5_addr; // @[SocTop.scala 27:32]
  assign io_sram5_cen = sram_bridge_io_sram_share_5_cen; // @[SocTop.scala 27:32]
  assign io_sram5_wen = sram_bridge_io_sram_share_5_wen; // @[SocTop.scala 27:32]
  assign io_sram5_wdata = sram_bridge_io_sram_share_5_wdata; // @[SocTop.scala 27:32]
  assign io_sram6_addr = sram_bridge_io_sram_share_6_addr; // @[SocTop.scala 28:32]
  assign io_sram6_cen = sram_bridge_io_sram_share_6_cen; // @[SocTop.scala 28:32]
  assign io_sram6_wen = sram_bridge_io_sram_share_6_wen; // @[SocTop.scala 28:32]
  assign io_sram6_wdata = sram_bridge_io_sram_share_6_wdata; // @[SocTop.scala 28:32]
  assign io_sram7_addr = sram_bridge_io_sram_share_7_addr; // @[SocTop.scala 29:32]
  assign io_sram7_cen = sram_bridge_io_sram_share_7_cen; // @[SocTop.scala 29:32]
  assign io_sram7_wen = sram_bridge_io_sram_share_7_wen; // @[SocTop.scala 29:32]
  assign io_sram7_wdata = sram_bridge_io_sram_share_7_wdata; // @[SocTop.scala 29:32]
  assign io_commit_0_pc = core_io_commit_0_pc;
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_icache_bridge_rd_rdy = transfer_bridge_io_icache_rd_rdy; // @[SocTop.scala 32:29]
  assign core_io_icache_bridge_ret_valid = transfer_bridge_io_icache_ret_valid; // @[SocTop.scala 32:29]
  assign core_io_icache_bridge_ret_data = transfer_bridge_io_icache_ret_data; // @[SocTop.scala 32:29]
  assign core_io_dcache_bridge_rd_rdy = transfer_bridge_io_dcache_rd_rdy; // @[SocTop.scala 33:29]
  assign core_io_dcache_bridge_ret_valid = transfer_bridge_io_dcache_ret_valid; // @[SocTop.scala 33:29]
  assign core_io_dcache_bridge_ret_data = transfer_bridge_io_dcache_ret_data; // @[SocTop.scala 33:29]
  assign core_io_dcache_bridge_wr_rdy = transfer_bridge_io_dcache_wr_rdy; // @[SocTop.scala 33:29]
  assign core_io_dcache_bridge_wr_ok = transfer_bridge_io_dcache_wr_ok; // @[SocTop.scala 33:29]
  assign core_io_sram_0_rdata = sram_bridge_io_sram_cache_0_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_1_rdata = sram_bridge_io_sram_cache_1_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_2_rdata = sram_bridge_io_sram_cache_2_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_3_rdata = sram_bridge_io_sram_cache_3_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_4_rdata = sram_bridge_io_sram_cache_4_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_5_rdata = sram_bridge_io_sram_cache_5_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_6_rdata = sram_bridge_io_sram_cache_6_rdata; // @[SocTop.scala 21:29]
  assign core_io_sram_7_rdata = sram_bridge_io_sram_cache_7_rdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_0_en = core_io_sram_0_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_0_wen = core_io_sram_0_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_0_addr = core_io_sram_0_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_0_wdata = core_io_sram_0_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_1_en = core_io_sram_1_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_1_wen = core_io_sram_1_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_1_addr = core_io_sram_1_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_1_wdata = core_io_sram_1_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_2_en = core_io_sram_2_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_2_wen = core_io_sram_2_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_2_addr = core_io_sram_2_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_2_wdata = core_io_sram_2_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_3_en = core_io_sram_3_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_3_wen = core_io_sram_3_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_3_addr = core_io_sram_3_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_3_wdata = core_io_sram_3_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_4_en = core_io_sram_4_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_4_wen = core_io_sram_4_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_4_addr = core_io_sram_4_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_4_wdata = core_io_sram_4_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_5_en = core_io_sram_5_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_5_wen = core_io_sram_5_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_5_addr = core_io_sram_5_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_5_wdata = core_io_sram_5_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_6_en = core_io_sram_6_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_6_wen = core_io_sram_6_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_6_addr = core_io_sram_6_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_6_wdata = core_io_sram_6_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_7_en = core_io_sram_7_en; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_7_wen = core_io_sram_7_wen; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_7_addr = core_io_sram_7_addr; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_cache_7_wdata = core_io_sram_7_wdata; // @[SocTop.scala 21:29]
  assign sram_bridge_io_sram_share_0_rdata = io_sram0_rdata; // @[SocTop.scala 22:32]
  assign sram_bridge_io_sram_share_1_rdata = io_sram1_rdata; // @[SocTop.scala 23:32]
  assign sram_bridge_io_sram_share_2_rdata = io_sram2_rdata; // @[SocTop.scala 24:32]
  assign sram_bridge_io_sram_share_3_rdata = io_sram3_rdata; // @[SocTop.scala 25:32]
  assign sram_bridge_io_sram_share_4_rdata = io_sram4_rdata; // @[SocTop.scala 26:32]
  assign sram_bridge_io_sram_share_5_rdata = io_sram5_rdata; // @[SocTop.scala 27:32]
  assign sram_bridge_io_sram_share_6_rdata = io_sram6_rdata; // @[SocTop.scala 28:32]
  assign sram_bridge_io_sram_share_7_rdata = io_sram7_rdata; // @[SocTop.scala 29:32]
  assign transfer_bridge_clock = clock;
  assign transfer_bridge_reset = reset;
  assign transfer_bridge_io_icache_rd_req = core_io_icache_bridge_rd_req; // @[SocTop.scala 32:29]
  assign transfer_bridge_io_icache_rd_size = core_io_icache_bridge_rd_size; // @[SocTop.scala 32:29]
  assign transfer_bridge_io_icache_rd_addr = core_io_icache_bridge_rd_addr; // @[SocTop.scala 32:29]
  assign transfer_bridge_io_dcache_rd_req = core_io_dcache_bridge_rd_req; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_rd_size = core_io_dcache_bridge_rd_size; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_rd_addr = core_io_dcache_bridge_rd_addr; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_wr_req = core_io_dcache_bridge_wr_req; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_wr_size = core_io_dcache_bridge_wr_size; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_wr_addr = core_io_dcache_bridge_wr_addr; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_wr_wstrb = core_io_dcache_bridge_wr_wstrb; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_dcache_wr_data = core_io_dcache_bridge_wr_data; // @[SocTop.scala 33:29]
  assign transfer_bridge_io_out_awready = io_master_awready; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_wready = io_master_wready; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_bvalid = io_master_bvalid; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_arready = io_master_arready; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_rvalid = io_master_rvalid; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_rdata = io_master_rdata; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_rlast = io_master_rlast; // @[SocTop.scala 34:26]
  assign transfer_bridge_io_out_rid = io_master_rid; // @[SocTop.scala 34:26]
endmodule
module SRAM(
  input          clock,
  input          io_en,
  input          io_wen,
  input  [5:0]   io_addr,
  input  [127:0] io_wdata,
  output [127:0] io_rdata
);
  wire [127:0] sram_Q; // @[SRAM.scala 52:20]
  wire  sram_CLK; // @[SRAM.scala 52:20]
  wire  sram_CEN; // @[SRAM.scala 52:20]
  wire  sram_WEN; // @[SRAM.scala 52:20]
  wire [5:0] sram_A; // @[SRAM.scala 52:20]
  wire [127:0] sram_D; // @[SRAM.scala 52:20]
  S011HD1P_X32Y2D128 sram ( // @[SRAM.scala 52:20]
    .Q(sram_Q),
    .CLK(sram_CLK),
    .CEN(sram_CEN),
    .WEN(sram_WEN),
    .A(sram_A),
    .D(sram_D)
  );
  assign io_rdata = sram_Q; // @[SRAM.scala 54:12]
  assign sram_CLK = clock; // @[SRAM.scala 56:15]
  assign sram_CEN = ~io_en; // @[SRAM.scala 57:18]
  assign sram_WEN = ~io_wen; // @[SRAM.scala 58:18]
  assign sram_A = io_addr; // @[SRAM.scala 59:13]
  assign sram_D = io_wdata; // @[SRAM.scala 60:13]
endmodule
module MySimTop(
  input         clock,
  input         reset,
  input         io_axi_awready,
  output        io_axi_awvalid,
  output [31:0] io_axi_awaddr,
  output [3:0]  io_axi_awid,
  output [7:0]  io_axi_awlen,
  output [2:0]  io_axi_awsize,
  output [1:0]  io_axi_awburst,
  input         io_axi_wready,
  output        io_axi_wvalid,
  output [63:0] io_axi_wdata,
  output [7:0]  io_axi_wstrb,
  output        io_axi_wlast,
  output        io_axi_bready,
  input         io_axi_bvalid,
  input  [1:0]  io_axi_bresp,
  input  [3:0]  io_axi_bid,
  input         io_axi_arready,
  output        io_axi_arvalid,
  output [31:0] io_axi_araddr,
  output [3:0]  io_axi_arid,
  output [7:0]  io_axi_arlen,
  output [2:0]  io_axi_arsize,
  output [1:0]  io_axi_arburst,
  output        io_axi_rready,
  input         io_axi_rvalid,
  input  [1:0]  io_axi_rresp,
  input  [63:0] io_axi_rdata,
  input         io_axi_rlast,
  input  [3:0]  io_axi_rid,
  output [31:0] io_pc
);
  wire  soctop_clock; // @[MySimTop.scala 12:22]
  wire  soctop_reset; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_awready; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_awvalid; // @[MySimTop.scala 12:22]
  wire [31:0] soctop_io_master_awaddr; // @[MySimTop.scala 12:22]
  wire [7:0] soctop_io_master_awlen; // @[MySimTop.scala 12:22]
  wire [2:0] soctop_io_master_awsize; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_wready; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_wvalid; // @[MySimTop.scala 12:22]
  wire [63:0] soctop_io_master_wdata; // @[MySimTop.scala 12:22]
  wire [7:0] soctop_io_master_wstrb; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_wlast; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_bready; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_bvalid; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_arready; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_arvalid; // @[MySimTop.scala 12:22]
  wire [31:0] soctop_io_master_araddr; // @[MySimTop.scala 12:22]
  wire [3:0] soctop_io_master_arid; // @[MySimTop.scala 12:22]
  wire [7:0] soctop_io_master_arlen; // @[MySimTop.scala 12:22]
  wire [2:0] soctop_io_master_arsize; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_rvalid; // @[MySimTop.scala 12:22]
  wire [63:0] soctop_io_master_rdata; // @[MySimTop.scala 12:22]
  wire  soctop_io_master_rlast; // @[MySimTop.scala 12:22]
  wire [3:0] soctop_io_master_rid; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram0_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram0_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram0_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram0_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram0_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram1_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram1_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram1_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram1_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram1_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram2_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram2_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram2_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram2_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram2_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram3_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram3_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram3_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram3_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram3_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram4_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram4_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram4_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram4_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram4_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram5_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram5_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram5_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram5_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram5_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram6_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram6_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram6_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram6_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram6_rdata; // @[MySimTop.scala 12:22]
  wire [5:0] soctop_io_sram7_addr; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram7_cen; // @[MySimTop.scala 12:22]
  wire  soctop_io_sram7_wen; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram7_wdata; // @[MySimTop.scala 12:22]
  wire [127:0] soctop_io_sram7_rdata; // @[MySimTop.scala 12:22]
  wire [31:0] soctop_io_commit_0_pc; // @[MySimTop.scala 12:22]
  wire  sram_0_clock; // @[MySimTop.scala 26:22]
  wire  sram_0_io_en; // @[MySimTop.scala 26:22]
  wire  sram_0_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_0_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_0_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_0_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_1_clock; // @[MySimTop.scala 26:22]
  wire  sram_1_io_en; // @[MySimTop.scala 26:22]
  wire  sram_1_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_1_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_1_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_1_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_2_clock; // @[MySimTop.scala 26:22]
  wire  sram_2_io_en; // @[MySimTop.scala 26:22]
  wire  sram_2_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_2_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_2_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_2_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_3_clock; // @[MySimTop.scala 26:22]
  wire  sram_3_io_en; // @[MySimTop.scala 26:22]
  wire  sram_3_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_3_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_3_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_3_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_4_clock; // @[MySimTop.scala 26:22]
  wire  sram_4_io_en; // @[MySimTop.scala 26:22]
  wire  sram_4_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_4_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_4_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_4_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_5_clock; // @[MySimTop.scala 26:22]
  wire  sram_5_io_en; // @[MySimTop.scala 26:22]
  wire  sram_5_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_5_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_5_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_5_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_6_clock; // @[MySimTop.scala 26:22]
  wire  sram_6_io_en; // @[MySimTop.scala 26:22]
  wire  sram_6_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_6_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_6_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_6_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_7_clock; // @[MySimTop.scala 26:22]
  wire  sram_7_io_en; // @[MySimTop.scala 26:22]
  wire  sram_7_io_wen; // @[MySimTop.scala 26:22]
  wire [5:0] sram_7_io_addr; // @[MySimTop.scala 26:22]
  wire [127:0] sram_7_io_wdata; // @[MySimTop.scala 26:22]
  wire [127:0] sram_7_io_rdata; // @[MySimTop.scala 26:22]
  wire  sram_from_soctop_0_cen = soctop_io_sram0_cen; // @[MySimTop.scala 15:30 MySimTop.scala 16:23]
  wire  sram_from_soctop_0_wen = soctop_io_sram0_wen; // @[MySimTop.scala 15:30 MySimTop.scala 16:23]
  wire  sram_from_soctop_1_cen = soctop_io_sram1_cen; // @[MySimTop.scala 15:30 MySimTop.scala 17:23]
  wire  sram_from_soctop_1_wen = soctop_io_sram1_wen; // @[MySimTop.scala 15:30 MySimTop.scala 17:23]
  wire  sram_from_soctop_2_cen = soctop_io_sram2_cen; // @[MySimTop.scala 15:30 MySimTop.scala 18:23]
  wire  sram_from_soctop_2_wen = soctop_io_sram2_wen; // @[MySimTop.scala 15:30 MySimTop.scala 18:23]
  wire  sram_from_soctop_3_cen = soctop_io_sram3_cen; // @[MySimTop.scala 15:30 MySimTop.scala 19:23]
  wire  sram_from_soctop_3_wen = soctop_io_sram3_wen; // @[MySimTop.scala 15:30 MySimTop.scala 19:23]
  wire  sram_from_soctop_4_cen = soctop_io_sram4_cen; // @[MySimTop.scala 15:30 MySimTop.scala 20:23]
  wire  sram_from_soctop_4_wen = soctop_io_sram4_wen; // @[MySimTop.scala 15:30 MySimTop.scala 20:23]
  wire  sram_from_soctop_5_cen = soctop_io_sram5_cen; // @[MySimTop.scala 15:30 MySimTop.scala 21:23]
  wire  sram_from_soctop_5_wen = soctop_io_sram5_wen; // @[MySimTop.scala 15:30 MySimTop.scala 21:23]
  wire  sram_from_soctop_6_cen = soctop_io_sram6_cen; // @[MySimTop.scala 15:30 MySimTop.scala 22:23]
  wire  sram_from_soctop_6_wen = soctop_io_sram6_wen; // @[MySimTop.scala 15:30 MySimTop.scala 22:23]
  wire  sram_from_soctop_7_cen = soctop_io_sram7_cen; // @[MySimTop.scala 15:30 MySimTop.scala 23:23]
  wire  sram_from_soctop_7_wen = soctop_io_sram7_wen; // @[MySimTop.scala 15:30 MySimTop.scala 23:23]
  SocTop soctop ( // @[MySimTop.scala 12:22]
    .clock(soctop_clock),
    .reset(soctop_reset),
    .io_master_awready(soctop_io_master_awready),
    .io_master_awvalid(soctop_io_master_awvalid),
    .io_master_awaddr(soctop_io_master_awaddr),
    .io_master_awlen(soctop_io_master_awlen),
    .io_master_awsize(soctop_io_master_awsize),
    .io_master_wready(soctop_io_master_wready),
    .io_master_wvalid(soctop_io_master_wvalid),
    .io_master_wdata(soctop_io_master_wdata),
    .io_master_wstrb(soctop_io_master_wstrb),
    .io_master_wlast(soctop_io_master_wlast),
    .io_master_bready(soctop_io_master_bready),
    .io_master_bvalid(soctop_io_master_bvalid),
    .io_master_arready(soctop_io_master_arready),
    .io_master_arvalid(soctop_io_master_arvalid),
    .io_master_araddr(soctop_io_master_araddr),
    .io_master_arid(soctop_io_master_arid),
    .io_master_arlen(soctop_io_master_arlen),
    .io_master_arsize(soctop_io_master_arsize),
    .io_master_rvalid(soctop_io_master_rvalid),
    .io_master_rdata(soctop_io_master_rdata),
    .io_master_rlast(soctop_io_master_rlast),
    .io_master_rid(soctop_io_master_rid),
    .io_sram0_addr(soctop_io_sram0_addr),
    .io_sram0_cen(soctop_io_sram0_cen),
    .io_sram0_wen(soctop_io_sram0_wen),
    .io_sram0_wdata(soctop_io_sram0_wdata),
    .io_sram0_rdata(soctop_io_sram0_rdata),
    .io_sram1_addr(soctop_io_sram1_addr),
    .io_sram1_cen(soctop_io_sram1_cen),
    .io_sram1_wen(soctop_io_sram1_wen),
    .io_sram1_wdata(soctop_io_sram1_wdata),
    .io_sram1_rdata(soctop_io_sram1_rdata),
    .io_sram2_addr(soctop_io_sram2_addr),
    .io_sram2_cen(soctop_io_sram2_cen),
    .io_sram2_wen(soctop_io_sram2_wen),
    .io_sram2_wdata(soctop_io_sram2_wdata),
    .io_sram2_rdata(soctop_io_sram2_rdata),
    .io_sram3_addr(soctop_io_sram3_addr),
    .io_sram3_cen(soctop_io_sram3_cen),
    .io_sram3_wen(soctop_io_sram3_wen),
    .io_sram3_wdata(soctop_io_sram3_wdata),
    .io_sram3_rdata(soctop_io_sram3_rdata),
    .io_sram4_addr(soctop_io_sram4_addr),
    .io_sram4_cen(soctop_io_sram4_cen),
    .io_sram4_wen(soctop_io_sram4_wen),
    .io_sram4_wdata(soctop_io_sram4_wdata),
    .io_sram4_rdata(soctop_io_sram4_rdata),
    .io_sram5_addr(soctop_io_sram5_addr),
    .io_sram5_cen(soctop_io_sram5_cen),
    .io_sram5_wen(soctop_io_sram5_wen),
    .io_sram5_wdata(soctop_io_sram5_wdata),
    .io_sram5_rdata(soctop_io_sram5_rdata),
    .io_sram6_addr(soctop_io_sram6_addr),
    .io_sram6_cen(soctop_io_sram6_cen),
    .io_sram6_wen(soctop_io_sram6_wen),
    .io_sram6_wdata(soctop_io_sram6_wdata),
    .io_sram6_rdata(soctop_io_sram6_rdata),
    .io_sram7_addr(soctop_io_sram7_addr),
    .io_sram7_cen(soctop_io_sram7_cen),
    .io_sram7_wen(soctop_io_sram7_wen),
    .io_sram7_wdata(soctop_io_sram7_wdata),
    .io_sram7_rdata(soctop_io_sram7_rdata),
    .io_commit_0_pc(soctop_io_commit_0_pc)
  );
  SRAM sram_0 ( // @[MySimTop.scala 26:22]
    .clock(sram_0_clock),
    .io_en(sram_0_io_en),
    .io_wen(sram_0_io_wen),
    .io_addr(sram_0_io_addr),
    .io_wdata(sram_0_io_wdata),
    .io_rdata(sram_0_io_rdata)
  );
  SRAM sram_1 ( // @[MySimTop.scala 26:22]
    .clock(sram_1_clock),
    .io_en(sram_1_io_en),
    .io_wen(sram_1_io_wen),
    .io_addr(sram_1_io_addr),
    .io_wdata(sram_1_io_wdata),
    .io_rdata(sram_1_io_rdata)
  );
  SRAM sram_2 ( // @[MySimTop.scala 26:22]
    .clock(sram_2_clock),
    .io_en(sram_2_io_en),
    .io_wen(sram_2_io_wen),
    .io_addr(sram_2_io_addr),
    .io_wdata(sram_2_io_wdata),
    .io_rdata(sram_2_io_rdata)
  );
  SRAM sram_3 ( // @[MySimTop.scala 26:22]
    .clock(sram_3_clock),
    .io_en(sram_3_io_en),
    .io_wen(sram_3_io_wen),
    .io_addr(sram_3_io_addr),
    .io_wdata(sram_3_io_wdata),
    .io_rdata(sram_3_io_rdata)
  );
  SRAM sram_4 ( // @[MySimTop.scala 26:22]
    .clock(sram_4_clock),
    .io_en(sram_4_io_en),
    .io_wen(sram_4_io_wen),
    .io_addr(sram_4_io_addr),
    .io_wdata(sram_4_io_wdata),
    .io_rdata(sram_4_io_rdata)
  );
  SRAM sram_5 ( // @[MySimTop.scala 26:22]
    .clock(sram_5_clock),
    .io_en(sram_5_io_en),
    .io_wen(sram_5_io_wen),
    .io_addr(sram_5_io_addr),
    .io_wdata(sram_5_io_wdata),
    .io_rdata(sram_5_io_rdata)
  );
  SRAM sram_6 ( // @[MySimTop.scala 26:22]
    .clock(sram_6_clock),
    .io_en(sram_6_io_en),
    .io_wen(sram_6_io_wen),
    .io_addr(sram_6_io_addr),
    .io_wdata(sram_6_io_wdata),
    .io_rdata(sram_6_io_rdata)
  );
  SRAM sram_7 ( // @[MySimTop.scala 26:22]
    .clock(sram_7_clock),
    .io_en(sram_7_io_en),
    .io_wen(sram_7_io_wen),
    .io_addr(sram_7_io_addr),
    .io_wdata(sram_7_io_wdata),
    .io_rdata(sram_7_io_rdata)
  );
  assign io_axi_awvalid = soctop_io_master_awvalid; // @[MySimTop.scala 13:10]
  assign io_axi_awaddr = soctop_io_master_awaddr; // @[MySimTop.scala 13:10]
  assign io_axi_awid = 4'h1; // @[MySimTop.scala 13:10]
  assign io_axi_awlen = soctop_io_master_awlen; // @[MySimTop.scala 13:10]
  assign io_axi_awsize = soctop_io_master_awsize; // @[MySimTop.scala 13:10]
  assign io_axi_awburst = 2'h1; // @[MySimTop.scala 13:10]
  assign io_axi_wvalid = soctop_io_master_wvalid; // @[MySimTop.scala 13:10]
  assign io_axi_wdata = soctop_io_master_wdata; // @[MySimTop.scala 13:10]
  assign io_axi_wstrb = soctop_io_master_wstrb; // @[MySimTop.scala 13:10]
  assign io_axi_wlast = soctop_io_master_wlast; // @[MySimTop.scala 13:10]
  assign io_axi_bready = soctop_io_master_bready; // @[MySimTop.scala 13:10]
  assign io_axi_arvalid = soctop_io_master_arvalid; // @[MySimTop.scala 13:10]
  assign io_axi_araddr = soctop_io_master_araddr; // @[MySimTop.scala 13:10]
  assign io_axi_arid = soctop_io_master_arid; // @[MySimTop.scala 13:10]
  assign io_axi_arlen = soctop_io_master_arlen; // @[MySimTop.scala 13:10]
  assign io_axi_arsize = soctop_io_master_arsize; // @[MySimTop.scala 13:10]
  assign io_axi_arburst = 2'h1; // @[MySimTop.scala 13:10]
  assign io_axi_rready = 1'h1; // @[MySimTop.scala 13:10]
  assign io_pc = soctop_io_commit_0_pc;
  assign soctop_clock = clock;
  assign soctop_reset = reset;
  assign soctop_io_master_awready = io_axi_awready; // @[MySimTop.scala 13:10]
  assign soctop_io_master_wready = io_axi_wready; // @[MySimTop.scala 13:10]
  assign soctop_io_master_bvalid = io_axi_bvalid; // @[MySimTop.scala 13:10]
  assign soctop_io_master_arready = io_axi_arready; // @[MySimTop.scala 13:10]
  assign soctop_io_master_rvalid = io_axi_rvalid; // @[MySimTop.scala 13:10]
  assign soctop_io_master_rdata = io_axi_rdata; // @[MySimTop.scala 13:10]
  assign soctop_io_master_rlast = io_axi_rlast; // @[MySimTop.scala 13:10]
  assign soctop_io_master_rid = io_axi_rid; // @[MySimTop.scala 13:10]
  assign soctop_io_sram0_rdata = sram_0_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram1_rdata = sram_1_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram2_rdata = sram_2_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram3_rdata = sram_3_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram4_rdata = sram_4_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram5_rdata = sram_5_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram6_rdata = sram_6_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign soctop_io_sram7_rdata = sram_7_io_rdata; // @[MySimTop.scala 15:30 MySimTop.scala 36:31]
  assign sram_0_clock = clock;
  assign sram_0_io_en = ~sram_from_soctop_0_cen; // @[MySimTop.scala 32:22]
  assign sram_0_io_wen = ~sram_from_soctop_0_wen; // @[MySimTop.scala 33:23]
  assign sram_0_io_addr = soctop_io_sram0_addr; // @[MySimTop.scala 15:30 MySimTop.scala 16:23]
  assign sram_0_io_wdata = soctop_io_sram0_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 16:23]
  assign sram_1_clock = clock;
  assign sram_1_io_en = ~sram_from_soctop_1_cen; // @[MySimTop.scala 32:22]
  assign sram_1_io_wen = ~sram_from_soctop_1_wen; // @[MySimTop.scala 33:23]
  assign sram_1_io_addr = soctop_io_sram1_addr; // @[MySimTop.scala 15:30 MySimTop.scala 17:23]
  assign sram_1_io_wdata = soctop_io_sram1_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 17:23]
  assign sram_2_clock = clock;
  assign sram_2_io_en = ~sram_from_soctop_2_cen; // @[MySimTop.scala 32:22]
  assign sram_2_io_wen = ~sram_from_soctop_2_wen; // @[MySimTop.scala 33:23]
  assign sram_2_io_addr = soctop_io_sram2_addr; // @[MySimTop.scala 15:30 MySimTop.scala 18:23]
  assign sram_2_io_wdata = soctop_io_sram2_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 18:23]
  assign sram_3_clock = clock;
  assign sram_3_io_en = ~sram_from_soctop_3_cen; // @[MySimTop.scala 32:22]
  assign sram_3_io_wen = ~sram_from_soctop_3_wen; // @[MySimTop.scala 33:23]
  assign sram_3_io_addr = soctop_io_sram3_addr; // @[MySimTop.scala 15:30 MySimTop.scala 19:23]
  assign sram_3_io_wdata = soctop_io_sram3_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 19:23]
  assign sram_4_clock = clock;
  assign sram_4_io_en = ~sram_from_soctop_4_cen; // @[MySimTop.scala 32:22]
  assign sram_4_io_wen = ~sram_from_soctop_4_wen; // @[MySimTop.scala 33:23]
  assign sram_4_io_addr = soctop_io_sram4_addr; // @[MySimTop.scala 15:30 MySimTop.scala 20:23]
  assign sram_4_io_wdata = soctop_io_sram4_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 20:23]
  assign sram_5_clock = clock;
  assign sram_5_io_en = ~sram_from_soctop_5_cen; // @[MySimTop.scala 32:22]
  assign sram_5_io_wen = ~sram_from_soctop_5_wen; // @[MySimTop.scala 33:23]
  assign sram_5_io_addr = soctop_io_sram5_addr; // @[MySimTop.scala 15:30 MySimTop.scala 21:23]
  assign sram_5_io_wdata = soctop_io_sram5_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 21:23]
  assign sram_6_clock = clock;
  assign sram_6_io_en = ~sram_from_soctop_6_cen; // @[MySimTop.scala 32:22]
  assign sram_6_io_wen = ~sram_from_soctop_6_wen; // @[MySimTop.scala 33:23]
  assign sram_6_io_addr = soctop_io_sram6_addr; // @[MySimTop.scala 15:30 MySimTop.scala 22:23]
  assign sram_6_io_wdata = soctop_io_sram6_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 22:23]
  assign sram_7_clock = clock;
  assign sram_7_io_en = ~sram_from_soctop_7_cen; // @[MySimTop.scala 32:22]
  assign sram_7_io_wen = ~sram_from_soctop_7_wen; // @[MySimTop.scala 33:23]
  assign sram_7_io_addr = soctop_io_sram7_addr; // @[MySimTop.scala 15:30 MySimTop.scala 23:23]
  assign sram_7_io_wdata = soctop_io_sram7_wdata; // @[MySimTop.scala 15:30 MySimTop.scala 23:23]
endmodule
